magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect 0 0 664 806
<< pmoslvt >>
rect 204 102 304 704
rect 360 102 460 704
<< pdiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 304 692 360 704
rect 304 658 315 692
rect 349 658 360 692
rect 304 624 360 658
rect 304 590 315 624
rect 349 590 360 624
rect 304 556 360 590
rect 304 522 315 556
rect 349 522 360 556
rect 304 488 360 522
rect 304 454 315 488
rect 349 454 360 488
rect 304 420 360 454
rect 304 386 315 420
rect 349 386 360 420
rect 304 352 360 386
rect 304 318 315 352
rect 349 318 360 352
rect 304 284 360 318
rect 304 250 315 284
rect 349 250 360 284
rect 304 216 360 250
rect 304 182 315 216
rect 349 182 360 216
rect 304 148 360 182
rect 304 114 315 148
rect 349 114 360 148
rect 304 102 360 114
rect 460 692 516 704
rect 460 658 471 692
rect 505 658 516 692
rect 460 624 516 658
rect 460 590 471 624
rect 505 590 516 624
rect 460 556 516 590
rect 460 522 471 556
rect 505 522 516 556
rect 460 488 516 522
rect 460 454 471 488
rect 505 454 516 488
rect 460 420 516 454
rect 460 386 471 420
rect 505 386 516 420
rect 460 352 516 386
rect 460 318 471 352
rect 505 318 516 352
rect 460 284 516 318
rect 460 250 471 284
rect 505 250 516 284
rect 460 216 516 250
rect 460 182 471 216
rect 505 182 516 216
rect 460 148 516 182
rect 460 114 471 148
rect 505 114 516 148
rect 460 102 516 114
<< pdiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 315 658 349 692
rect 315 590 349 624
rect 315 522 349 556
rect 315 454 349 488
rect 315 386 349 420
rect 315 318 349 352
rect 315 250 349 284
rect 315 182 349 216
rect 315 114 349 148
rect 471 658 505 692
rect 471 590 505 624
rect 471 522 505 556
rect 471 454 505 488
rect 471 386 505 420
rect 471 318 505 352
rect 471 250 505 284
rect 471 182 505 216
rect 471 114 505 148
<< nsubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 570 658 628 704
rect 570 624 582 658
rect 616 624 628 658
rect 570 590 628 624
rect 570 556 582 590
rect 616 556 628 590
rect 570 522 628 556
rect 570 488 582 522
rect 616 488 628 522
rect 570 454 628 488
rect 570 420 582 454
rect 616 420 628 454
rect 570 386 628 420
rect 570 352 582 386
rect 616 352 628 386
rect 570 318 628 352
rect 570 284 582 318
rect 616 284 628 318
rect 570 250 628 284
rect 570 216 582 250
rect 616 216 628 250
rect 570 182 628 216
rect 570 148 582 182
rect 616 148 628 182
rect 570 102 628 148
<< nsubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 582 624 616 658
rect 582 556 616 590
rect 582 488 616 522
rect 582 420 616 454
rect 582 352 616 386
rect 582 284 616 318
rect 582 216 616 250
rect 582 148 616 182
<< poly >>
rect 159 786 505 806
rect 159 752 179 786
rect 213 752 247 786
rect 281 752 315 786
rect 349 752 383 786
rect 417 752 451 786
rect 485 752 505 786
rect 159 736 505 752
rect 204 704 304 736
rect 360 704 460 736
rect 204 70 304 102
rect 360 70 460 102
rect 159 54 505 70
rect 159 20 179 54
rect 213 20 247 54
rect 281 20 315 54
rect 349 20 383 54
rect 417 20 451 54
rect 485 20 505 54
rect 159 0 505 20
<< polycont >>
rect 179 752 213 786
rect 247 752 281 786
rect 315 752 349 786
rect 383 752 417 786
rect 451 752 485 786
rect 179 20 213 54
rect 247 20 281 54
rect 315 20 349 54
rect 383 20 417 54
rect 451 20 485 54
<< locali >>
rect 159 752 171 786
rect 213 752 243 786
rect 281 752 315 786
rect 349 752 383 786
rect 421 752 451 786
rect 493 752 505 786
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 315 692 349 708
rect 315 624 349 638
rect 315 556 349 566
rect 315 488 349 494
rect 315 420 349 422
rect 315 384 349 386
rect 315 312 349 318
rect 315 240 349 250
rect 315 168 349 182
rect 315 98 349 114
rect 471 692 505 708
rect 471 624 505 638
rect 471 556 505 566
rect 471 488 505 494
rect 471 420 505 422
rect 471 384 505 386
rect 471 312 505 318
rect 471 240 505 250
rect 471 168 505 182
rect 582 672 616 674
rect 582 600 616 624
rect 582 528 616 556
rect 582 456 616 488
rect 582 386 616 420
rect 582 318 616 350
rect 582 250 616 278
rect 582 182 616 206
rect 582 132 616 134
rect 471 98 505 114
rect 159 20 171 54
rect 213 20 243 54
rect 281 20 315 54
rect 349 20 383 54
rect 421 20 451 54
rect 493 20 505 54
<< viali >>
rect 171 752 179 786
rect 179 752 205 786
rect 243 752 247 786
rect 247 752 277 786
rect 315 752 349 786
rect 387 752 417 786
rect 417 752 421 786
rect 459 752 485 786
rect 485 752 493 786
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 315 658 349 672
rect 315 638 349 658
rect 315 590 349 600
rect 315 566 349 590
rect 315 522 349 528
rect 315 494 349 522
rect 315 454 349 456
rect 315 422 349 454
rect 315 352 349 384
rect 315 350 349 352
rect 315 284 349 312
rect 315 278 349 284
rect 315 216 349 240
rect 315 206 349 216
rect 315 148 349 168
rect 315 134 349 148
rect 471 658 505 672
rect 471 638 505 658
rect 471 590 505 600
rect 471 566 505 590
rect 471 522 505 528
rect 471 494 505 522
rect 471 454 505 456
rect 471 422 505 454
rect 471 352 505 384
rect 471 350 505 352
rect 471 284 505 312
rect 471 278 505 284
rect 471 216 505 240
rect 471 206 505 216
rect 471 148 505 168
rect 471 134 505 148
rect 582 658 616 672
rect 582 638 616 658
rect 582 590 616 600
rect 582 566 616 590
rect 582 522 616 528
rect 582 494 616 522
rect 582 454 616 456
rect 582 422 616 454
rect 582 352 616 384
rect 582 350 616 352
rect 582 284 616 312
rect 582 278 616 284
rect 582 216 616 240
rect 582 206 616 216
rect 582 148 616 168
rect 582 134 616 148
rect 171 20 179 54
rect 179 20 205 54
rect 243 20 247 54
rect 247 20 277 54
rect 315 20 349 54
rect 387 20 417 54
rect 417 20 421 54
rect 459 20 485 54
rect 485 20 493 54
<< metal1 >>
rect 159 786 505 806
rect 159 752 171 786
rect 205 752 243 786
rect 277 752 315 786
rect 349 752 387 786
rect 421 752 459 786
rect 493 752 505 786
rect 159 740 505 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 306 678 358 684
rect 306 614 358 626
rect 306 550 358 562
rect 306 494 315 498
rect 349 494 358 498
rect 306 486 358 494
rect 306 422 315 434
rect 349 422 358 434
rect 306 384 358 422
rect 306 350 315 384
rect 349 350 358 384
rect 306 312 358 350
rect 306 278 315 312
rect 349 278 358 312
rect 306 240 358 278
rect 306 206 315 240
rect 349 206 358 240
rect 306 168 358 206
rect 306 134 315 168
rect 349 134 358 168
rect 306 122 358 134
rect 462 672 514 684
rect 462 638 471 672
rect 505 638 514 672
rect 462 600 514 638
rect 462 566 471 600
rect 505 566 514 600
rect 462 528 514 566
rect 462 494 471 528
rect 505 494 514 528
rect 462 456 514 494
rect 462 422 471 456
rect 505 422 514 456
rect 462 384 514 422
rect 462 372 471 384
rect 505 372 514 384
rect 462 312 514 320
rect 462 308 471 312
rect 505 308 514 312
rect 462 244 514 256
rect 462 180 514 192
rect 462 122 514 128
rect 570 672 628 684
rect 570 638 582 672
rect 616 638 628 672
rect 570 600 628 638
rect 570 566 582 600
rect 616 566 628 600
rect 570 528 628 566
rect 570 494 582 528
rect 616 494 628 528
rect 570 456 628 494
rect 570 422 582 456
rect 616 422 628 456
rect 570 384 628 422
rect 570 350 582 384
rect 616 350 628 384
rect 570 312 628 350
rect 570 278 582 312
rect 616 278 628 312
rect 570 240 628 278
rect 570 206 582 240
rect 616 206 628 240
rect 570 168 628 206
rect 570 134 582 168
rect 616 134 628 168
rect 570 122 628 134
rect 159 54 505 66
rect 159 20 171 54
rect 205 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 505 54
rect 159 0 505 20
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 306 672 358 678
rect 306 638 315 672
rect 315 638 349 672
rect 349 638 358 672
rect 306 626 358 638
rect 306 600 358 614
rect 306 566 315 600
rect 315 566 349 600
rect 349 566 358 600
rect 306 562 358 566
rect 306 528 358 550
rect 306 498 315 528
rect 315 498 349 528
rect 349 498 358 528
rect 306 456 358 486
rect 306 434 315 456
rect 315 434 349 456
rect 349 434 358 456
rect 462 350 471 372
rect 471 350 505 372
rect 505 350 514 372
rect 462 320 514 350
rect 462 278 471 308
rect 471 278 505 308
rect 505 278 514 308
rect 462 256 514 278
rect 462 240 514 244
rect 462 206 471 240
rect 471 206 505 240
rect 505 206 514 240
rect 462 192 514 206
rect 462 168 514 180
rect 462 134 471 168
rect 471 134 505 168
rect 505 134 514 168
rect 462 128 514 134
<< metal2 >>
rect 10 678 654 684
rect 10 626 306 678
rect 358 626 654 678
rect 10 614 654 626
rect 10 562 306 614
rect 358 562 654 614
rect 10 550 654 562
rect 10 498 306 550
rect 358 498 654 550
rect 10 486 654 498
rect 10 434 306 486
rect 358 434 654 486
rect 10 428 654 434
rect 10 372 654 378
rect 10 320 150 372
rect 202 320 462 372
rect 514 320 654 372
rect 10 308 654 320
rect 10 256 150 308
rect 202 256 462 308
rect 514 256 654 308
rect 10 244 654 256
rect 10 192 150 244
rect 202 192 462 244
rect 514 192 654 244
rect 10 180 654 192
rect 10 128 150 180
rect 202 128 462 180
rect 514 128 654 180
rect 10 122 654 128
<< labels >>
flabel metal2 s 10 122 30 378 7 FreeSans 300 180 0 0 SOURCE
flabel metal2 s 10 428 30 684 7 FreeSans 300 180 0 0 DRAIN
flabel metal1 s 159 740 505 806 0 FreeSans 300 0 0 0 GATE
flabel metal1 s 159 0 505 66 0 FreeSans 300 0 0 0 GATE
flabel metal1 s 570 122 628 138 3 FreeSans 300 90 0 0 BULK
flabel metal1 s 36 122 94 138 3 FreeSans 300 90 0 0 BULK
<< properties >>
string GDS_END 9979256
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9967764
<< end >>
