/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice