/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hvl/lef/sky130_fd_sc_hvl.lef