magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< locali >>
rect 7840 50423 7899 50457
rect 11965 50423 11993 50457
rect 7865 50278 7899 50423
rect 7865 50244 7958 50278
rect 7865 50052 7958 50086
rect 7865 49907 7899 50052
rect 7840 49873 7899 49907
rect 11965 49873 11993 49907
rect 7840 49633 7899 49667
rect 11965 49633 11993 49667
rect 7865 49488 7899 49633
rect 7865 49454 7958 49488
rect 7865 49262 7958 49296
rect 7865 49117 7899 49262
rect 7840 49083 7899 49117
rect 11965 49083 11993 49117
rect 7840 48843 7899 48877
rect 11965 48843 11993 48877
rect 7865 48698 7899 48843
rect 7865 48664 7958 48698
rect 7865 48472 7958 48506
rect 7865 48327 7899 48472
rect 7840 48293 7899 48327
rect 11965 48293 11993 48327
rect 7840 48053 7899 48087
rect 11965 48053 11993 48087
rect 7865 47908 7899 48053
rect 7865 47874 7958 47908
rect 7865 47682 7958 47716
rect 7865 47537 7899 47682
rect 7840 47503 7899 47537
rect 11965 47503 11993 47537
rect 7840 47263 7899 47297
rect 11965 47263 11993 47297
rect 7865 47118 7899 47263
rect 7865 47084 7958 47118
rect 7865 46892 7958 46926
rect 7865 46747 7899 46892
rect 7840 46713 7899 46747
rect 11965 46713 11993 46747
rect 7840 46473 7899 46507
rect 11965 46473 11993 46507
rect 7865 46328 7899 46473
rect 7865 46294 7958 46328
rect 7865 46102 7958 46136
rect 7865 45957 7899 46102
rect 7840 45923 7899 45957
rect 11965 45923 11993 45957
rect 7840 45683 7899 45717
rect 11965 45683 11993 45717
rect 7865 45538 7899 45683
rect 7865 45504 7958 45538
rect 7865 45312 7958 45346
rect 7865 45167 7899 45312
rect 7840 45133 7899 45167
rect 11965 45133 11993 45167
rect 7840 44893 7899 44927
rect 11965 44893 11993 44927
rect 7865 44748 7899 44893
rect 7865 44714 7958 44748
rect 7865 44522 7958 44556
rect 7865 44377 7899 44522
rect 7840 44343 7899 44377
rect 11965 44343 11993 44377
rect 7840 44103 7899 44137
rect 11965 44103 11993 44137
rect 7865 43958 7899 44103
rect 7865 43924 7958 43958
rect 7865 43732 7958 43766
rect 7865 43587 7899 43732
rect 7840 43553 7899 43587
rect 11965 43553 11993 43587
rect 7840 43313 7899 43347
rect 11965 43313 11993 43347
rect 7865 43168 7899 43313
rect 7865 43134 7958 43168
rect 7865 42942 7958 42976
rect 7865 42797 7899 42942
rect 7840 42763 7899 42797
rect 11965 42763 11993 42797
rect 7840 42523 7899 42557
rect 11965 42523 11993 42557
rect 7865 42378 7899 42523
rect 7865 42344 7958 42378
rect 7865 42152 7958 42186
rect 7865 42007 7899 42152
rect 7840 41973 7899 42007
rect 11965 41973 11993 42007
rect 7840 41733 7899 41767
rect 11965 41733 11993 41767
rect 7865 41588 7899 41733
rect 7865 41554 7958 41588
rect 7865 41362 7958 41396
rect 7865 41217 7899 41362
rect 7840 41183 7899 41217
rect 11965 41183 11993 41217
rect 7840 40943 7899 40977
rect 11965 40943 11993 40977
rect 7865 40798 7899 40943
rect 7865 40764 7958 40798
rect 7865 40572 7958 40606
rect 7865 40427 7899 40572
rect 7840 40393 7899 40427
rect 11965 40393 11993 40427
rect 7840 40153 7899 40187
rect 11965 40153 11993 40187
rect 7865 40008 7899 40153
rect 7865 39974 7958 40008
rect 7865 39782 7958 39816
rect 7865 39637 7899 39782
rect 7840 39603 7899 39637
rect 11965 39603 11993 39637
rect 7840 39363 7899 39397
rect 11965 39363 11993 39397
rect 7865 39218 7899 39363
rect 7865 39184 7958 39218
rect 7865 38992 7958 39026
rect 7865 38847 7899 38992
rect 7840 38813 7899 38847
rect 11965 38813 11993 38847
rect 7840 38573 7899 38607
rect 11965 38573 11993 38607
rect 7865 38428 7899 38573
rect 7865 38394 7958 38428
rect 7865 38202 7958 38236
rect 7865 38057 7899 38202
rect 7840 38023 7899 38057
rect 11965 38023 11993 38057
rect 7840 37783 7899 37817
rect 11965 37783 11993 37817
rect 7865 37638 7899 37783
rect 7865 37604 7958 37638
rect 7865 37412 7958 37446
rect 7865 37267 7899 37412
rect 7840 37233 7899 37267
rect 11965 37233 11993 37267
rect 7840 36993 7899 37027
rect 11965 36993 11993 37027
rect 7865 36848 7899 36993
rect 7865 36814 7958 36848
rect 7865 36622 7958 36656
rect 7865 36477 7899 36622
rect 7840 36443 7899 36477
rect 11965 36443 11993 36477
rect 7840 36203 7899 36237
rect 11965 36203 11993 36237
rect 7865 36058 7899 36203
rect 7865 36024 7958 36058
rect 7865 35832 7958 35866
rect 7865 35687 7899 35832
rect 7840 35653 7899 35687
rect 11965 35653 11993 35687
rect 7840 35413 7899 35447
rect 11965 35413 11993 35447
rect 7865 35268 7899 35413
rect 7865 35234 7958 35268
rect 7865 35042 7958 35076
rect 7865 34897 7899 35042
rect 7840 34863 7899 34897
rect 11965 34863 11993 34897
rect 7840 34623 7899 34657
rect 11965 34623 11993 34657
rect 7865 34478 7899 34623
rect 7865 34444 7958 34478
rect 7865 34252 7958 34286
rect 7865 34107 7899 34252
rect 7840 34073 7899 34107
rect 11965 34073 11993 34107
rect 7840 33833 7899 33867
rect 11965 33833 11993 33867
rect 7865 33688 7899 33833
rect 7865 33654 7958 33688
rect 7865 33462 7958 33496
rect 7865 33317 7899 33462
rect 7840 33283 7899 33317
rect 11965 33283 11993 33317
rect 7840 33043 7899 33077
rect 11965 33043 11993 33077
rect 7865 32898 7899 33043
rect 7865 32864 7958 32898
rect 7865 32672 7958 32706
rect 7865 32527 7899 32672
rect 7840 32493 7899 32527
rect 11965 32493 11993 32527
rect 7840 32253 7899 32287
rect 11965 32253 11993 32287
rect 7865 32108 7899 32253
rect 7865 32074 7958 32108
rect 7865 31882 7958 31916
rect 7865 31737 7899 31882
rect 7840 31703 7899 31737
rect 11965 31703 11993 31737
rect 7840 31463 7899 31497
rect 11965 31463 11993 31497
rect 7865 31318 7899 31463
rect 7865 31284 7958 31318
rect 7865 31092 7958 31126
rect 7865 30947 7899 31092
rect 7840 30913 7899 30947
rect 11965 30913 11993 30947
rect 7840 30673 7899 30707
rect 11965 30673 11993 30707
rect 7865 30528 7899 30673
rect 7865 30494 7958 30528
rect 7865 30302 7958 30336
rect 7865 30157 7899 30302
rect 7840 30123 7899 30157
rect 11965 30123 11993 30157
rect 7840 29883 7899 29917
rect 11965 29883 11993 29917
rect 7865 29738 7899 29883
rect 7865 29704 7958 29738
rect 7865 29512 7958 29546
rect 7865 29367 7899 29512
rect 7840 29333 7899 29367
rect 11965 29333 11993 29367
rect 7840 29093 7899 29127
rect 11965 29093 11993 29127
rect 7865 28948 7899 29093
rect 7865 28914 7958 28948
rect 7865 28722 7958 28756
rect 7865 28577 7899 28722
rect 7840 28543 7899 28577
rect 11965 28543 11993 28577
rect 7840 28303 7899 28337
rect 11965 28303 11993 28337
rect 7865 28158 7899 28303
rect 7865 28124 7958 28158
rect 7865 27932 7958 27966
rect 7865 27787 7899 27932
rect 7840 27753 7899 27787
rect 11965 27753 11993 27787
rect 7840 27513 7899 27547
rect 11965 27513 11993 27547
rect 7865 27368 7899 27513
rect 7865 27334 7958 27368
rect 7865 27142 7958 27176
rect 7865 26997 7899 27142
rect 7840 26963 7899 26997
rect 11965 26963 11993 26997
rect 7840 26723 7899 26757
rect 11965 26723 11993 26757
rect 7865 26578 7899 26723
rect 7865 26544 7958 26578
rect 7865 26352 7958 26386
rect 7865 26207 7899 26352
rect 7840 26173 7899 26207
rect 11965 26173 11993 26207
rect 7840 25933 7899 25967
rect 11965 25933 11993 25967
rect 7865 25788 7899 25933
rect 7865 25754 7958 25788
rect 7865 25562 7958 25596
rect 7865 25417 7899 25562
rect 7840 25383 7899 25417
rect 11965 25383 11993 25417
rect 7840 25143 7899 25177
rect 11965 25143 11993 25177
rect 7865 24998 7899 25143
rect 7865 24964 7958 24998
rect 7865 24772 7958 24806
rect 7865 24627 7899 24772
rect 7840 24593 7899 24627
rect 11965 24593 11993 24627
rect 7840 24353 7899 24387
rect 11965 24353 11993 24387
rect 7865 24208 7899 24353
rect 7865 24174 7958 24208
rect 7865 23982 7958 24016
rect 7865 23837 7899 23982
rect 7840 23803 7899 23837
rect 11965 23803 11993 23837
rect 7840 23563 7899 23597
rect 11965 23563 11993 23597
rect 7865 23418 7899 23563
rect 7865 23384 7958 23418
rect 7865 23192 7958 23226
rect 7865 23047 7899 23192
rect 7840 23013 7899 23047
rect 11965 23013 11993 23047
rect 7840 22773 7899 22807
rect 11965 22773 11993 22807
rect 7865 22628 7899 22773
rect 7865 22594 7958 22628
rect 7865 22402 7958 22436
rect 7865 22257 7899 22402
rect 7840 22223 7899 22257
rect 11965 22223 11993 22257
rect 7840 21983 7899 22017
rect 11965 21983 11993 22017
rect 7865 21838 7899 21983
rect 7865 21804 7958 21838
rect 7865 21612 7958 21646
rect 7865 21467 7899 21612
rect 7840 21433 7899 21467
rect 11965 21433 11993 21467
rect 7840 21193 7899 21227
rect 11965 21193 11993 21227
rect 7865 21048 7899 21193
rect 7865 21014 7958 21048
rect 7865 20822 7958 20856
rect 7865 20677 7899 20822
rect 7840 20643 7899 20677
rect 11965 20643 11993 20677
rect 7840 20403 7899 20437
rect 11965 20403 11993 20437
rect 7865 20258 7899 20403
rect 7865 20224 7958 20258
rect 7865 20032 7958 20066
rect 7865 19887 7899 20032
rect 7840 19853 7899 19887
rect 11965 19853 11993 19887
rect 7840 19613 7899 19647
rect 11965 19613 11993 19647
rect 7865 19468 7899 19613
rect 7865 19434 7958 19468
rect 7865 19242 7958 19276
rect 7865 19097 7899 19242
rect 7840 19063 7899 19097
rect 11965 19063 11993 19097
rect 7840 18823 7899 18857
rect 11965 18823 11993 18857
rect 7865 18678 7899 18823
rect 7865 18644 7958 18678
rect 7865 18452 7958 18486
rect 7865 18307 7899 18452
rect 7840 18273 7899 18307
rect 11965 18273 11993 18307
rect 7840 18033 7899 18067
rect 11965 18033 11993 18067
rect 7865 17888 7899 18033
rect 7865 17854 7958 17888
rect 7865 17662 7958 17696
rect 7865 17517 7899 17662
rect 7840 17483 7899 17517
rect 11965 17483 11993 17517
rect 7840 17243 7899 17277
rect 11965 17243 11993 17277
rect 7865 17098 7899 17243
rect 7865 17064 7958 17098
rect 7865 16872 7958 16906
rect 7865 16727 7899 16872
rect 7840 16693 7899 16727
rect 11965 16693 11993 16727
rect 7840 16453 7899 16487
rect 11965 16453 11993 16487
rect 7865 16308 7899 16453
rect 7865 16274 7958 16308
rect 7865 16082 7958 16116
rect 7865 15937 7899 16082
rect 7840 15903 7899 15937
rect 11965 15903 11993 15937
rect 7840 15663 7899 15697
rect 11965 15663 11993 15697
rect 7865 15518 7899 15663
rect 7865 15484 7958 15518
rect 7865 15292 7958 15326
rect 7865 15147 7899 15292
rect 7840 15113 7899 15147
rect 11965 15113 11993 15147
rect 7840 14873 7899 14907
rect 11965 14873 11993 14907
rect 7865 14728 7899 14873
rect 7865 14694 7958 14728
rect 7865 14502 7958 14536
rect 7865 14357 7899 14502
rect 7840 14323 7899 14357
rect 11965 14323 11993 14357
rect 7840 14083 7899 14117
rect 11965 14083 11993 14117
rect 7865 13938 7899 14083
rect 7865 13904 7958 13938
rect 7865 13712 7958 13746
rect 7865 13567 7899 13712
rect 7840 13533 7899 13567
rect 11965 13533 11993 13567
rect 7840 13293 7899 13327
rect 11965 13293 11993 13327
rect 7865 13148 7899 13293
rect 7865 13114 7958 13148
rect 7865 12922 7958 12956
rect 7865 12777 7899 12922
rect 7840 12743 7899 12777
rect 11965 12743 11993 12777
rect 7840 12503 7899 12537
rect 11965 12503 11993 12537
rect 7865 12358 7899 12503
rect 7865 12324 7958 12358
rect 7865 12132 7958 12166
rect 7865 11987 7899 12132
rect 7840 11953 7899 11987
rect 11965 11953 11993 11987
rect 7840 11713 7899 11747
rect 11965 11713 11993 11747
rect 7865 11568 7899 11713
rect 7865 11534 7958 11568
rect 7865 11342 7958 11376
rect 7865 11197 7899 11342
rect 7840 11163 7899 11197
rect 11965 11163 11993 11197
rect 7840 10923 7899 10957
rect 11965 10923 11993 10957
rect 7865 10778 7899 10923
rect 7865 10744 7958 10778
rect 7865 10552 7958 10586
rect 7865 10407 7899 10552
rect 7840 10373 7899 10407
rect 11965 10373 11993 10407
rect 7840 10133 7899 10167
rect 11965 10133 11993 10167
rect 7865 9988 7899 10133
rect 7865 9954 7958 9988
rect 7865 9762 7958 9796
rect 7865 9617 7899 9762
rect 7840 9583 7899 9617
rect 11965 9583 11993 9617
rect 7840 9343 7899 9377
rect 11965 9343 11993 9377
rect 7865 9198 7899 9343
rect 7865 9164 7958 9198
rect 7865 8972 7958 9006
rect 7865 8827 7899 8972
rect 7840 8793 7899 8827
rect 11965 8793 11993 8827
rect 7840 8553 7899 8587
rect 11965 8553 11993 8587
rect 7865 8408 7899 8553
rect 7865 8374 7958 8408
rect 7865 8182 7958 8216
rect 7865 8037 7899 8182
rect 7840 8003 7899 8037
rect 11965 8003 11993 8037
rect 7840 7763 7899 7797
rect 11965 7763 11993 7797
rect 7865 7618 7899 7763
rect 7865 7584 7958 7618
rect 7865 7392 7958 7426
rect 7865 7247 7899 7392
rect 7840 7213 7899 7247
rect 11965 7213 11993 7247
rect 7840 6973 7899 7007
rect 11965 6973 11993 7007
rect 7865 6828 7899 6973
rect 7865 6794 7958 6828
rect 7865 6602 7958 6636
rect 7865 6457 7899 6602
rect 7840 6423 7899 6457
rect 11965 6423 11993 6457
rect 7840 6183 7899 6217
rect 11965 6183 11993 6217
rect 7865 6038 7899 6183
rect 7865 6004 7958 6038
rect 7865 5812 7958 5846
rect 7865 5667 7899 5812
rect 7840 5633 7899 5667
rect 11965 5633 11993 5667
rect 7840 5393 7899 5427
rect 11965 5393 11993 5427
rect 7865 5248 7899 5393
rect 7865 5214 7958 5248
rect 7865 5022 7958 5056
rect 7865 4877 7899 5022
rect 7840 4843 7899 4877
rect 11965 4843 11993 4877
rect 7840 4603 7899 4637
rect 11965 4603 11993 4637
rect 7865 4458 7899 4603
rect 7865 4424 7958 4458
rect 7865 4232 7958 4266
rect 7865 4087 7899 4232
rect 7840 4053 7899 4087
rect 11965 4053 11993 4087
rect 7840 3813 7899 3847
rect 11965 3813 11993 3847
rect 7865 3668 7899 3813
rect 7865 3634 7958 3668
rect 7865 3442 7958 3476
rect 7865 3297 7899 3442
rect 7840 3263 7899 3297
rect 11965 3263 11993 3297
rect 7840 3023 7899 3057
rect 11965 3023 11993 3057
rect 7865 2878 7899 3023
rect 7865 2844 7958 2878
rect 7865 2652 7958 2686
rect 7865 2507 7899 2652
rect 7840 2473 7899 2507
rect 11965 2473 11993 2507
rect 7840 2233 7899 2267
rect 11965 2233 11993 2267
rect 7865 2088 7899 2233
rect 7865 2054 7958 2088
rect 7865 1862 7958 1896
rect 7865 1717 7899 1862
rect 7840 1683 7899 1717
rect 11965 1683 11993 1717
rect 7840 1443 7899 1477
rect 11965 1443 11993 1477
rect 7865 1298 7899 1443
rect 7865 1264 7958 1298
rect 7865 1072 7958 1106
rect 7865 927 7899 1072
rect 7840 893 7899 927
rect 11965 893 11993 927
rect 7840 653 7899 687
rect 11965 653 11993 687
rect 7865 508 7899 653
rect 7865 474 7958 508
rect 7865 282 7958 316
rect 7865 137 7899 282
rect 7840 103 7899 137
rect 11965 103 11993 137
rect 9576 -137 11993 -103
rect 7717 -174 7751 -158
rect 7751 -208 7974 -174
rect 7717 -224 7751 -208
rect 7957 -282 7991 -266
rect 7957 -332 7991 -316
<< viali >>
rect 7717 -208 7751 -174
rect 7957 -316 7991 -282
<< metal1 >>
rect 8109 25239 8115 25291
rect 8167 25239 8173 25291
rect 8534 25238 8540 25290
rect 8592 25238 8598 25290
rect 9577 25254 9583 25306
rect 9635 25254 9641 25306
rect 11225 25254 11231 25306
rect 11283 25254 11289 25306
rect 19 0 47 7900
rect 99 0 127 7900
rect 179 0 207 7900
rect 259 0 287 7900
rect 339 0 367 7900
rect 419 0 447 7900
rect 499 0 527 7900
rect 7702 -217 7708 -165
rect 7760 -217 7766 -165
rect 8534 -211 8540 -159
rect 8592 -211 8598 -159
rect 11225 -224 11231 -172
rect 11283 -224 11289 -172
rect 7942 -325 7948 -273
rect 8000 -325 8006 -273
<< via1 >>
rect 8115 25239 8167 25291
rect 8540 25238 8592 25290
rect 9583 25254 9635 25306
rect 11231 25254 11283 25306
rect 7708 -174 7760 -165
rect 7708 -208 7717 -174
rect 7717 -208 7751 -174
rect 7751 -208 7760 -174
rect 7708 -217 7760 -208
rect 8540 -211 8592 -159
rect 11231 -224 11283 -172
rect 7948 -282 8000 -273
rect 7948 -316 7957 -282
rect 7957 -316 7991 -282
rect 7991 -316 8000 -282
rect 7948 -325 8000 -316
<< metal2 >>
rect 9581 25308 9637 25317
rect 8113 25293 8169 25302
rect 8113 25228 8169 25237
rect 8538 25292 8594 25301
rect 9581 25243 9637 25252
rect 11229 25308 11285 25317
rect 11229 25243 11285 25252
rect 8538 25227 8594 25236
rect 7941 -136 7969 0
rect 7706 -163 7762 -154
rect 7941 -164 7988 -136
rect 7706 -228 7762 -219
rect 7960 -267 7988 -164
rect 8538 -157 8594 -148
rect 8538 -222 8594 -213
rect 11229 -169 11285 -160
rect 11229 -234 11285 -225
rect 7948 -273 8000 -267
rect 7948 -331 8000 -325
<< via2 >>
rect 9581 25306 9637 25308
rect 8113 25291 8169 25293
rect 8113 25239 8115 25291
rect 8115 25239 8167 25291
rect 8167 25239 8169 25291
rect 8113 25237 8169 25239
rect 8538 25290 8594 25292
rect 8538 25238 8540 25290
rect 8540 25238 8592 25290
rect 8592 25238 8594 25290
rect 9581 25254 9583 25306
rect 9583 25254 9635 25306
rect 9635 25254 9637 25306
rect 9581 25252 9637 25254
rect 11229 25306 11285 25308
rect 11229 25254 11231 25306
rect 11231 25254 11283 25306
rect 11283 25254 11285 25306
rect 11229 25252 11285 25254
rect 8538 25236 8594 25238
rect 7706 -165 7762 -163
rect 7706 -217 7708 -165
rect 7708 -217 7760 -165
rect 7760 -217 7762 -165
rect 7706 -219 7762 -217
rect 8538 -159 8594 -157
rect 8538 -211 8540 -159
rect 8540 -211 8592 -159
rect 8592 -211 8594 -159
rect 8538 -213 8594 -211
rect 11229 -172 11285 -169
rect 11229 -224 11231 -172
rect 11231 -224 11283 -172
rect 11283 -224 11285 -172
rect 11229 -225 11285 -224
<< metal3 >>
rect 6025 50139 6123 50237
rect 6450 50139 6548 50237
rect 6882 50139 6980 50237
rect 7264 50116 7362 50214
rect 7660 50116 7758 50214
rect 6025 49765 6123 49863
rect 6450 49707 6548 49805
rect 6882 49707 6980 49805
rect 7264 49721 7362 49819
rect 7660 49721 7758 49819
rect 6025 49349 6123 49447
rect 6450 49349 6548 49447
rect 6882 49349 6980 49447
rect 7264 49326 7362 49424
rect 7660 49326 7758 49424
rect 6025 48975 6123 49073
rect 6450 48917 6548 49015
rect 6882 48917 6980 49015
rect 7264 48931 7362 49029
rect 7660 48931 7758 49029
rect 6025 48559 6123 48657
rect 6450 48559 6548 48657
rect 6882 48559 6980 48657
rect 7264 48536 7362 48634
rect 7660 48536 7758 48634
rect 6025 48185 6123 48283
rect 6450 48127 6548 48225
rect 6882 48127 6980 48225
rect 7264 48141 7362 48239
rect 7660 48141 7758 48239
rect 6025 47769 6123 47867
rect 6450 47769 6548 47867
rect 6882 47769 6980 47867
rect 7264 47746 7362 47844
rect 7660 47746 7758 47844
rect 6025 47395 6123 47493
rect 6450 47337 6548 47435
rect 6882 47337 6980 47435
rect 7264 47351 7362 47449
rect 7660 47351 7758 47449
rect 6025 46979 6123 47077
rect 6450 46979 6548 47077
rect 6882 46979 6980 47077
rect 7264 46956 7362 47054
rect 7660 46956 7758 47054
rect 6025 46605 6123 46703
rect 6450 46547 6548 46645
rect 6882 46547 6980 46645
rect 7264 46561 7362 46659
rect 7660 46561 7758 46659
rect 6025 46189 6123 46287
rect 6450 46189 6548 46287
rect 6882 46189 6980 46287
rect 7264 46166 7362 46264
rect 7660 46166 7758 46264
rect 6025 45815 6123 45913
rect 6450 45757 6548 45855
rect 6882 45757 6980 45855
rect 7264 45771 7362 45869
rect 7660 45771 7758 45869
rect 6025 45399 6123 45497
rect 6450 45399 6548 45497
rect 6882 45399 6980 45497
rect 7264 45376 7362 45474
rect 7660 45376 7758 45474
rect 6025 45025 6123 45123
rect 6450 44967 6548 45065
rect 6882 44967 6980 45065
rect 7264 44981 7362 45079
rect 7660 44981 7758 45079
rect 6025 44609 6123 44707
rect 6450 44609 6548 44707
rect 6882 44609 6980 44707
rect 7264 44586 7362 44684
rect 7660 44586 7758 44684
rect 6025 44235 6123 44333
rect 6450 44177 6548 44275
rect 6882 44177 6980 44275
rect 7264 44191 7362 44289
rect 7660 44191 7758 44289
rect 6025 43819 6123 43917
rect 6450 43819 6548 43917
rect 6882 43819 6980 43917
rect 7264 43796 7362 43894
rect 7660 43796 7758 43894
rect 6025 43445 6123 43543
rect 6450 43387 6548 43485
rect 6882 43387 6980 43485
rect 7264 43401 7362 43499
rect 7660 43401 7758 43499
rect 6025 43029 6123 43127
rect 6450 43029 6548 43127
rect 6882 43029 6980 43127
rect 7264 43006 7362 43104
rect 7660 43006 7758 43104
rect 6025 42655 6123 42753
rect 6450 42597 6548 42695
rect 6882 42597 6980 42695
rect 7264 42611 7362 42709
rect 7660 42611 7758 42709
rect 6025 42239 6123 42337
rect 6450 42239 6548 42337
rect 6882 42239 6980 42337
rect 7264 42216 7362 42314
rect 7660 42216 7758 42314
rect 6025 41865 6123 41963
rect 6450 41807 6548 41905
rect 6882 41807 6980 41905
rect 7264 41821 7362 41919
rect 7660 41821 7758 41919
rect 6025 41449 6123 41547
rect 6450 41449 6548 41547
rect 6882 41449 6980 41547
rect 7264 41426 7362 41524
rect 7660 41426 7758 41524
rect 6025 41075 6123 41173
rect 6450 41017 6548 41115
rect 6882 41017 6980 41115
rect 7264 41031 7362 41129
rect 7660 41031 7758 41129
rect 6025 40659 6123 40757
rect 6450 40659 6548 40757
rect 6882 40659 6980 40757
rect 7264 40636 7362 40734
rect 7660 40636 7758 40734
rect 6025 40285 6123 40383
rect 6450 40227 6548 40325
rect 6882 40227 6980 40325
rect 7264 40241 7362 40339
rect 7660 40241 7758 40339
rect 6025 39869 6123 39967
rect 6450 39869 6548 39967
rect 6882 39869 6980 39967
rect 7264 39846 7362 39944
rect 7660 39846 7758 39944
rect 6025 39495 6123 39593
rect 6450 39437 6548 39535
rect 6882 39437 6980 39535
rect 7264 39451 7362 39549
rect 7660 39451 7758 39549
rect 6025 39079 6123 39177
rect 6450 39079 6548 39177
rect 6882 39079 6980 39177
rect 7264 39056 7362 39154
rect 7660 39056 7758 39154
rect 6025 38705 6123 38803
rect 6450 38647 6548 38745
rect 6882 38647 6980 38745
rect 7264 38661 7362 38759
rect 7660 38661 7758 38759
rect 6025 38289 6123 38387
rect 6450 38289 6548 38387
rect 6882 38289 6980 38387
rect 7264 38266 7362 38364
rect 7660 38266 7758 38364
rect 6025 37915 6123 38013
rect 6450 37857 6548 37955
rect 6882 37857 6980 37955
rect 7264 37871 7362 37969
rect 7660 37871 7758 37969
rect 6025 37499 6123 37597
rect 6450 37499 6548 37597
rect 6882 37499 6980 37597
rect 7264 37476 7362 37574
rect 7660 37476 7758 37574
rect 6025 37125 6123 37223
rect 6450 37067 6548 37165
rect 6882 37067 6980 37165
rect 7264 37081 7362 37179
rect 7660 37081 7758 37179
rect 6025 36709 6123 36807
rect 6450 36709 6548 36807
rect 6882 36709 6980 36807
rect 7264 36686 7362 36784
rect 7660 36686 7758 36784
rect 6025 36335 6123 36433
rect 6450 36277 6548 36375
rect 6882 36277 6980 36375
rect 7264 36291 7362 36389
rect 7660 36291 7758 36389
rect 6025 35919 6123 36017
rect 6450 35919 6548 36017
rect 6882 35919 6980 36017
rect 7264 35896 7362 35994
rect 7660 35896 7758 35994
rect 6025 35545 6123 35643
rect 6450 35487 6548 35585
rect 6882 35487 6980 35585
rect 7264 35501 7362 35599
rect 7660 35501 7758 35599
rect 6025 35129 6123 35227
rect 6450 35129 6548 35227
rect 6882 35129 6980 35227
rect 7264 35106 7362 35204
rect 7660 35106 7758 35204
rect 6025 34755 6123 34853
rect 6450 34697 6548 34795
rect 6882 34697 6980 34795
rect 7264 34711 7362 34809
rect 7660 34711 7758 34809
rect 6025 34339 6123 34437
rect 6450 34339 6548 34437
rect 6882 34339 6980 34437
rect 7264 34316 7362 34414
rect 7660 34316 7758 34414
rect 6025 33965 6123 34063
rect 6450 33907 6548 34005
rect 6882 33907 6980 34005
rect 7264 33921 7362 34019
rect 7660 33921 7758 34019
rect 6025 33549 6123 33647
rect 6450 33549 6548 33647
rect 6882 33549 6980 33647
rect 7264 33526 7362 33624
rect 7660 33526 7758 33624
rect 6025 33175 6123 33273
rect 6450 33117 6548 33215
rect 6882 33117 6980 33215
rect 7264 33131 7362 33229
rect 7660 33131 7758 33229
rect 6025 32759 6123 32857
rect 6450 32759 6548 32857
rect 6882 32759 6980 32857
rect 7264 32736 7362 32834
rect 7660 32736 7758 32834
rect 6025 32385 6123 32483
rect 6450 32327 6548 32425
rect 6882 32327 6980 32425
rect 7264 32341 7362 32439
rect 7660 32341 7758 32439
rect 6025 31969 6123 32067
rect 6450 31969 6548 32067
rect 6882 31969 6980 32067
rect 7264 31946 7362 32044
rect 7660 31946 7758 32044
rect 6025 31595 6123 31693
rect 6450 31537 6548 31635
rect 6882 31537 6980 31635
rect 7264 31551 7362 31649
rect 7660 31551 7758 31649
rect 6025 31179 6123 31277
rect 6450 31179 6548 31277
rect 6882 31179 6980 31277
rect 7264 31156 7362 31254
rect 7660 31156 7758 31254
rect 6025 30805 6123 30903
rect 6450 30747 6548 30845
rect 6882 30747 6980 30845
rect 7264 30761 7362 30859
rect 7660 30761 7758 30859
rect 6025 30389 6123 30487
rect 6450 30389 6548 30487
rect 6882 30389 6980 30487
rect 7264 30366 7362 30464
rect 7660 30366 7758 30464
rect 6025 30015 6123 30113
rect 6450 29957 6548 30055
rect 6882 29957 6980 30055
rect 7264 29971 7362 30069
rect 7660 29971 7758 30069
rect 6025 29599 6123 29697
rect 6450 29599 6548 29697
rect 6882 29599 6980 29697
rect 7264 29576 7362 29674
rect 7660 29576 7758 29674
rect 6025 29225 6123 29323
rect 6450 29167 6548 29265
rect 6882 29167 6980 29265
rect 7264 29181 7362 29279
rect 7660 29181 7758 29279
rect 6025 28809 6123 28907
rect 6450 28809 6548 28907
rect 6882 28809 6980 28907
rect 7264 28786 7362 28884
rect 7660 28786 7758 28884
rect 6025 28435 6123 28533
rect 6450 28377 6548 28475
rect 6882 28377 6980 28475
rect 7264 28391 7362 28489
rect 7660 28391 7758 28489
rect 6025 28019 6123 28117
rect 6450 28019 6548 28117
rect 6882 28019 6980 28117
rect 7264 27996 7362 28094
rect 7660 27996 7758 28094
rect 6025 27645 6123 27743
rect 6450 27587 6548 27685
rect 6882 27587 6980 27685
rect 7264 27601 7362 27699
rect 7660 27601 7758 27699
rect 6025 27229 6123 27327
rect 6450 27229 6548 27327
rect 6882 27229 6980 27327
rect 7264 27206 7362 27304
rect 7660 27206 7758 27304
rect 6025 26855 6123 26953
rect 6450 26797 6548 26895
rect 6882 26797 6980 26895
rect 7264 26811 7362 26909
rect 7660 26811 7758 26909
rect 6025 26439 6123 26537
rect 6450 26439 6548 26537
rect 6882 26439 6980 26537
rect 7264 26416 7362 26514
rect 7660 26416 7758 26514
rect 6025 26065 6123 26163
rect 6450 26007 6548 26105
rect 6882 26007 6980 26105
rect 7264 26021 7362 26119
rect 7660 26021 7758 26119
rect 6025 25649 6123 25747
rect 6450 25649 6548 25747
rect 6882 25649 6980 25747
rect 7264 25626 7362 25724
rect 7660 25626 7758 25724
rect 6025 25275 6123 25373
rect 6450 25217 6548 25315
rect 6882 25217 6980 25315
rect 7264 25231 7362 25329
rect 7660 25231 7758 25329
rect 8092 25293 8190 25314
rect 8092 25237 8113 25293
rect 8169 25237 8190 25293
rect 8092 25216 8190 25237
rect 8517 25292 8615 25313
rect 8517 25236 8538 25292
rect 8594 25236 8615 25292
rect 8517 25215 8615 25236
rect 9560 25308 9658 25329
rect 9560 25252 9581 25308
rect 9637 25252 9658 25308
rect 9560 25231 9658 25252
rect 11208 25308 11306 25329
rect 11208 25252 11229 25308
rect 11285 25252 11306 25308
rect 11208 25231 11306 25252
rect 6025 24859 6123 24957
rect 6450 24859 6548 24957
rect 6882 24859 6980 24957
rect 7264 24836 7362 24934
rect 7660 24836 7758 24934
rect 6025 24485 6123 24583
rect 6450 24427 6548 24525
rect 6882 24427 6980 24525
rect 7264 24441 7362 24539
rect 7660 24441 7758 24539
rect 6025 24069 6123 24167
rect 6450 24069 6548 24167
rect 6882 24069 6980 24167
rect 7264 24046 7362 24144
rect 7660 24046 7758 24144
rect 6025 23695 6123 23793
rect 6450 23637 6548 23735
rect 6882 23637 6980 23735
rect 7264 23651 7362 23749
rect 7660 23651 7758 23749
rect 6025 23279 6123 23377
rect 6450 23279 6548 23377
rect 6882 23279 6980 23377
rect 7264 23256 7362 23354
rect 7660 23256 7758 23354
rect 6025 22905 6123 23003
rect 6450 22847 6548 22945
rect 6882 22847 6980 22945
rect 7264 22861 7362 22959
rect 7660 22861 7758 22959
rect 6025 22489 6123 22587
rect 6450 22489 6548 22587
rect 6882 22489 6980 22587
rect 7264 22466 7362 22564
rect 7660 22466 7758 22564
rect 6025 22115 6123 22213
rect 6450 22057 6548 22155
rect 6882 22057 6980 22155
rect 7264 22071 7362 22169
rect 7660 22071 7758 22169
rect 6025 21699 6123 21797
rect 6450 21699 6548 21797
rect 6882 21699 6980 21797
rect 7264 21676 7362 21774
rect 7660 21676 7758 21774
rect 6025 21325 6123 21423
rect 6450 21267 6548 21365
rect 6882 21267 6980 21365
rect 7264 21281 7362 21379
rect 7660 21281 7758 21379
rect 6025 20909 6123 21007
rect 6450 20909 6548 21007
rect 6882 20909 6980 21007
rect 7264 20886 7362 20984
rect 7660 20886 7758 20984
rect 6025 20535 6123 20633
rect 6450 20477 6548 20575
rect 6882 20477 6980 20575
rect 7264 20491 7362 20589
rect 7660 20491 7758 20589
rect 6025 20119 6123 20217
rect 6450 20119 6548 20217
rect 6882 20119 6980 20217
rect 7264 20096 7362 20194
rect 7660 20096 7758 20194
rect 6025 19745 6123 19843
rect 6450 19687 6548 19785
rect 6882 19687 6980 19785
rect 7264 19701 7362 19799
rect 7660 19701 7758 19799
rect 6025 19329 6123 19427
rect 6450 19329 6548 19427
rect 6882 19329 6980 19427
rect 7264 19306 7362 19404
rect 7660 19306 7758 19404
rect 6025 18955 6123 19053
rect 6450 18897 6548 18995
rect 6882 18897 6980 18995
rect 7264 18911 7362 19009
rect 7660 18911 7758 19009
rect 6025 18539 6123 18637
rect 6450 18539 6548 18637
rect 6882 18539 6980 18637
rect 7264 18516 7362 18614
rect 7660 18516 7758 18614
rect 6025 18165 6123 18263
rect 6450 18107 6548 18205
rect 6882 18107 6980 18205
rect 7264 18121 7362 18219
rect 7660 18121 7758 18219
rect 6025 17749 6123 17847
rect 6450 17749 6548 17847
rect 6882 17749 6980 17847
rect 7264 17726 7362 17824
rect 7660 17726 7758 17824
rect 6025 17375 6123 17473
rect 6450 17317 6548 17415
rect 6882 17317 6980 17415
rect 7264 17331 7362 17429
rect 7660 17331 7758 17429
rect 6025 16959 6123 17057
rect 6450 16959 6548 17057
rect 6882 16959 6980 17057
rect 7264 16936 7362 17034
rect 7660 16936 7758 17034
rect 6025 16585 6123 16683
rect 6450 16527 6548 16625
rect 6882 16527 6980 16625
rect 7264 16541 7362 16639
rect 7660 16541 7758 16639
rect 6025 16169 6123 16267
rect 6450 16169 6548 16267
rect 6882 16169 6980 16267
rect 7264 16146 7362 16244
rect 7660 16146 7758 16244
rect 6025 15795 6123 15893
rect 6450 15737 6548 15835
rect 6882 15737 6980 15835
rect 7264 15751 7362 15849
rect 7660 15751 7758 15849
rect 6025 15379 6123 15477
rect 6450 15379 6548 15477
rect 6882 15379 6980 15477
rect 7264 15356 7362 15454
rect 7660 15356 7758 15454
rect 6025 15005 6123 15103
rect 6450 14947 6548 15045
rect 6882 14947 6980 15045
rect 7264 14961 7362 15059
rect 7660 14961 7758 15059
rect 6025 14589 6123 14687
rect 6450 14589 6548 14687
rect 6882 14589 6980 14687
rect 7264 14566 7362 14664
rect 7660 14566 7758 14664
rect 6025 14215 6123 14313
rect 6450 14157 6548 14255
rect 6882 14157 6980 14255
rect 7264 14171 7362 14269
rect 7660 14171 7758 14269
rect 6025 13799 6123 13897
rect 6450 13799 6548 13897
rect 6882 13799 6980 13897
rect 7264 13776 7362 13874
rect 7660 13776 7758 13874
rect 6025 13425 6123 13523
rect 6450 13367 6548 13465
rect 6882 13367 6980 13465
rect 7264 13381 7362 13479
rect 7660 13381 7758 13479
rect 6025 13009 6123 13107
rect 6450 13009 6548 13107
rect 6882 13009 6980 13107
rect 7264 12986 7362 13084
rect 7660 12986 7758 13084
rect 6025 12635 6123 12733
rect 6450 12577 6548 12675
rect 6882 12577 6980 12675
rect 7264 12591 7362 12689
rect 7660 12591 7758 12689
rect 6025 12219 6123 12317
rect 6450 12219 6548 12317
rect 6882 12219 6980 12317
rect 7264 12196 7362 12294
rect 7660 12196 7758 12294
rect 6025 11845 6123 11943
rect 6450 11787 6548 11885
rect 6882 11787 6980 11885
rect 7264 11801 7362 11899
rect 7660 11801 7758 11899
rect 6025 11429 6123 11527
rect 6450 11429 6548 11527
rect 6882 11429 6980 11527
rect 7264 11406 7362 11504
rect 7660 11406 7758 11504
rect 6025 11055 6123 11153
rect 6450 10997 6548 11095
rect 6882 10997 6980 11095
rect 7264 11011 7362 11109
rect 7660 11011 7758 11109
rect 6025 10639 6123 10737
rect 6450 10639 6548 10737
rect 6882 10639 6980 10737
rect 7264 10616 7362 10714
rect 7660 10616 7758 10714
rect 6025 10265 6123 10363
rect 6450 10207 6548 10305
rect 6882 10207 6980 10305
rect 7264 10221 7362 10319
rect 7660 10221 7758 10319
rect 6025 9849 6123 9947
rect 6450 9849 6548 9947
rect 6882 9849 6980 9947
rect 7264 9826 7362 9924
rect 7660 9826 7758 9924
rect 6025 9475 6123 9573
rect 6450 9417 6548 9515
rect 6882 9417 6980 9515
rect 7264 9431 7362 9529
rect 7660 9431 7758 9529
rect 6025 9059 6123 9157
rect 6450 9059 6548 9157
rect 6882 9059 6980 9157
rect 7264 9036 7362 9134
rect 7660 9036 7758 9134
rect 6025 8685 6123 8783
rect 6450 8627 6548 8725
rect 6882 8627 6980 8725
rect 7264 8641 7362 8739
rect 7660 8641 7758 8739
rect 6025 8269 6123 8367
rect 6450 8269 6548 8367
rect 6882 8269 6980 8367
rect 7264 8246 7362 8344
rect 7660 8246 7758 8344
rect 6025 7895 6123 7993
rect 6450 7837 6548 7935
rect 6882 7837 6980 7935
rect 7264 7851 7362 7949
rect 7660 7851 7758 7949
rect 2611 7479 2709 7577
rect 3036 7479 3134 7577
rect 3468 7479 3566 7577
rect 3850 7456 3948 7554
rect 4246 7456 4344 7554
rect 6025 7479 6123 7577
rect 6450 7479 6548 7577
rect 6882 7479 6980 7577
rect 7264 7456 7362 7554
rect 7660 7456 7758 7554
rect 6025 7105 6123 7203
rect 6450 7047 6548 7145
rect 6882 7047 6980 7145
rect 7264 7061 7362 7159
rect 7660 7061 7758 7159
rect 2611 6689 2709 6787
rect 3036 6689 3134 6787
rect 3468 6689 3566 6787
rect 3850 6666 3948 6764
rect 4246 6666 4344 6764
rect 6025 6689 6123 6787
rect 6450 6689 6548 6787
rect 6882 6689 6980 6787
rect 7264 6666 7362 6764
rect 7660 6666 7758 6764
rect 6025 6315 6123 6413
rect 6450 6257 6548 6355
rect 6882 6257 6980 6355
rect 7264 6271 7362 6369
rect 7660 6271 7758 6369
rect 2611 5899 2709 5997
rect 3036 5899 3134 5997
rect 3468 5899 3566 5997
rect 3850 5876 3948 5974
rect 4246 5876 4344 5974
rect 6025 5899 6123 5997
rect 6450 5899 6548 5997
rect 6882 5899 6980 5997
rect 7264 5876 7362 5974
rect 7660 5876 7758 5974
rect 6025 5525 6123 5623
rect 6450 5467 6548 5565
rect 6882 5467 6980 5565
rect 7264 5481 7362 5579
rect 7660 5481 7758 5579
rect 1156 5086 1254 5184
rect 1552 5086 1650 5184
rect 2611 5109 2709 5207
rect 3036 5109 3134 5207
rect 3468 5109 3566 5207
rect 3850 5086 3948 5184
rect 4246 5086 4344 5184
rect 6025 5109 6123 5207
rect 6450 5109 6548 5207
rect 6882 5109 6980 5207
rect 7264 5086 7362 5184
rect 7660 5086 7758 5184
rect 6025 4735 6123 4833
rect 6450 4677 6548 4775
rect 6882 4677 6980 4775
rect 7264 4691 7362 4789
rect 7660 4691 7758 4789
rect 6025 4319 6123 4417
rect 6450 4319 6548 4417
rect 6882 4319 6980 4417
rect 7264 4296 7362 4394
rect 7660 4296 7758 4394
rect 6025 3945 6123 4043
rect 6450 3887 6548 3985
rect 6882 3887 6980 3985
rect 7264 3901 7362 3999
rect 7660 3901 7758 3999
rect 3046 3513 3144 3611
rect 3471 3513 3569 3611
rect 3850 3506 3948 3604
rect 4246 3506 4344 3604
rect 6025 3529 6123 3627
rect 6450 3529 6548 3627
rect 6882 3529 6980 3627
rect 7264 3506 7362 3604
rect 7660 3506 7758 3604
rect 6025 3155 6123 3253
rect 6450 3097 6548 3195
rect 6882 3097 6980 3195
rect 7264 3111 7362 3209
rect 7660 3111 7758 3209
rect 1752 2716 1850 2814
rect 2148 2716 2246 2814
rect 3046 2723 3144 2821
rect 3471 2723 3569 2821
rect 3850 2716 3948 2814
rect 4246 2716 4344 2814
rect 6025 2739 6123 2837
rect 6450 2739 6548 2837
rect 6882 2739 6980 2837
rect 7264 2716 7362 2814
rect 7660 2716 7758 2814
rect 6025 2365 6123 2463
rect 6450 2307 6548 2405
rect 6882 2307 6980 2405
rect 7264 2321 7362 2419
rect 7660 2321 7758 2419
rect 6025 1949 6123 2047
rect 6450 1949 6548 2047
rect 6882 1949 6980 2047
rect 7264 1926 7362 2024
rect 7660 1926 7758 2024
rect 6025 1575 6123 1673
rect 6450 1517 6548 1615
rect 6882 1517 6980 1615
rect 7264 1531 7362 1629
rect 7660 1531 7758 1629
rect 3046 1143 3144 1241
rect 3471 1143 3569 1241
rect 3850 1136 3948 1234
rect 4246 1136 4344 1234
rect 6025 1159 6123 1257
rect 6450 1159 6548 1257
rect 6882 1159 6980 1257
rect 7264 1136 7362 1234
rect 7660 1136 7758 1234
rect 6025 785 6123 883
rect 6450 727 6548 825
rect 6882 727 6980 825
rect 7264 741 7362 839
rect 7660 741 7758 839
rect 1752 346 1850 444
rect 2148 346 2246 444
rect 3046 353 3144 451
rect 3471 353 3569 451
rect 3850 346 3948 444
rect 4246 346 4344 444
rect 6025 369 6123 467
rect 6450 369 6548 467
rect 6882 369 6980 467
rect 7264 346 7362 444
rect 7660 346 7758 444
rect 7685 -163 7783 -142
rect 7685 -219 7706 -163
rect 7762 -219 7783 -163
rect 7685 -240 7783 -219
rect 8517 -157 8615 -136
rect 8517 -213 8538 -157
rect 8594 -213 8615 -157
rect 8517 -234 8615 -213
rect 11208 -169 11306 -148
rect 11208 -225 11229 -169
rect 11285 -225 11306 -169
rect 11208 -246 11306 -225
use sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_0  sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_0_0
timestamp 1676037725
transform 1 0 7871 0 -1 0
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_0
timestamp 1676037725
transform 1 0 7701 0 1 -228
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_1
timestamp 1676037725
transform 1 0 8533 0 1 -222
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_2
timestamp 1676037725
transform 1 0 11224 0 1 -234
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_3
timestamp 1676037725
transform 1 0 8108 0 1 25228
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_4
timestamp 1676037725
transform 1 0 9576 0 1 25243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_5
timestamp 1676037725
transform 1 0 8533 0 1 25227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_6
timestamp 1676037725
transform 1 0 11224 0 1 25243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_0
timestamp 1676037725
transform 1 0 7705 0 1 -224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_1
timestamp 1676037725
transform 1 0 7945 0 1 -332
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1676037725
transform 1 0 7702 0 1 -223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1676037725
transform 1 0 8534 0 1 -217
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1676037725
transform 1 0 11225 0 1 -230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_3
timestamp 1676037725
transform 1 0 8109 0 1 25233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_4
timestamp 1676037725
transform 1 0 9577 0 1 25248
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_5
timestamp 1676037725
transform 1 0 8534 0 1 25232
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_6
timestamp 1676037725
transform 1 0 11225 0 1 25248
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_7
timestamp 1676037725
transform 1 0 7942 0 1 -331
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder  sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0
timestamp 1676037725
transform 1 0 0 0 1 0
box 0 -60 7875 50620
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0
timestamp 1676037725
transform 1 0 7871 0 1 0
box 70 -56 4140 50616
<< labels >>
rlabel metal3 s 7660 48536 7758 48634 4 vdd
rlabel metal3 s 6450 46547 6548 46645 4 vdd
rlabel metal3 s 7660 45771 7758 45869 4 vdd
rlabel metal3 s 6882 46189 6980 46287 4 vdd
rlabel metal3 s 6882 46547 6980 46645 4 vdd
rlabel metal3 s 6450 48559 6548 48657 4 vdd
rlabel metal3 s 6450 46979 6548 47077 4 vdd
rlabel metal3 s 7660 49326 7758 49424 4 vdd
rlabel metal3 s 7660 46166 7758 46264 4 vdd
rlabel metal3 s 7660 44981 7758 45079 4 vdd
rlabel metal3 s 6882 45757 6980 45855 4 vdd
rlabel metal3 s 6450 44967 6548 45065 4 vdd
rlabel metal3 s 7660 50116 7758 50214 4 vdd
rlabel metal3 s 6882 47769 6980 47867 4 vdd
rlabel metal3 s 6882 44609 6980 44707 4 vdd
rlabel metal3 s 6450 50139 6548 50237 4 vdd
rlabel metal3 s 6450 44177 6548 44275 4 vdd
rlabel metal3 s 7660 47351 7758 47449 4 vdd
rlabel metal3 s 6450 45757 6548 45855 4 vdd
rlabel metal3 s 6450 47337 6548 47435 4 vdd
rlabel metal3 s 7660 49721 7758 49819 4 vdd
rlabel metal3 s 6450 49707 6548 49805 4 vdd
rlabel metal3 s 6882 44177 6980 44275 4 vdd
rlabel metal3 s 6450 48127 6548 48225 4 vdd
rlabel metal3 s 6882 47337 6980 47435 4 vdd
rlabel metal3 s 7660 48931 7758 49029 4 vdd
rlabel metal3 s 6882 48917 6980 49015 4 vdd
rlabel metal3 s 6450 48917 6548 49015 4 vdd
rlabel metal3 s 7660 48141 7758 48239 4 vdd
rlabel metal3 s 6882 44967 6980 45065 4 vdd
rlabel metal3 s 6882 49349 6980 49447 4 vdd
rlabel metal3 s 6882 45399 6980 45497 4 vdd
rlabel metal3 s 6882 46979 6980 47077 4 vdd
rlabel metal3 s 7660 46561 7758 46659 4 vdd
rlabel metal3 s 6882 49707 6980 49805 4 vdd
rlabel metal3 s 7660 47746 7758 47844 4 vdd
rlabel metal3 s 7660 46956 7758 47054 4 vdd
rlabel metal3 s 7660 44586 7758 44684 4 vdd
rlabel metal3 s 6450 49349 6548 49447 4 vdd
rlabel metal3 s 6450 44609 6548 44707 4 vdd
rlabel metal3 s 7660 45376 7758 45474 4 vdd
rlabel metal3 s 6882 48559 6980 48657 4 vdd
rlabel metal3 s 6450 46189 6548 46287 4 vdd
rlabel metal3 s 6450 45399 6548 45497 4 vdd
rlabel metal3 s 6882 50139 6980 50237 4 vdd
rlabel metal3 s 6882 48127 6980 48225 4 vdd
rlabel metal3 s 6450 47769 6548 47867 4 vdd
rlabel metal3 s 7660 44191 7758 44289 4 vdd
rlabel metal3 s 7264 44586 7362 44684 4 gnd
rlabel metal3 s 7264 45376 7362 45474 4 gnd
rlabel metal3 s 7264 46166 7362 46264 4 gnd
rlabel metal3 s 7264 47351 7362 47449 4 gnd
rlabel metal3 s 7264 48536 7362 48634 4 gnd
rlabel metal3 s 7264 47746 7362 47844 4 gnd
rlabel metal3 s 7264 44981 7362 45079 4 gnd
rlabel metal3 s 7264 48931 7362 49029 4 gnd
rlabel metal3 s 7264 49326 7362 49424 4 gnd
rlabel metal3 s 7264 46956 7362 47054 4 gnd
rlabel metal3 s 7264 44191 7362 44289 4 gnd
rlabel metal3 s 7264 50116 7362 50214 4 gnd
rlabel metal3 s 7264 48141 7362 48239 4 gnd
rlabel metal3 s 7264 45771 7362 45869 4 gnd
rlabel metal3 s 7264 46561 7362 46659 4 gnd
rlabel metal3 s 7264 49721 7362 49819 4 gnd
rlabel metal3 s 7660 38661 7758 38759 4 vdd
rlabel metal3 s 7660 41031 7758 41129 4 vdd
rlabel metal3 s 6450 39437 6548 39535 4 vdd
rlabel metal3 s 7660 37871 7758 37969 4 vdd
rlabel metal3 s 6450 43819 6548 43917 4 vdd
rlabel metal3 s 7660 43006 7758 43104 4 vdd
rlabel metal3 s 6882 41807 6980 41905 4 vdd
rlabel metal3 s 7660 42611 7758 42709 4 vdd
rlabel metal3 s 7660 39846 7758 39944 4 vdd
rlabel metal3 s 6450 40227 6548 40325 4 vdd
rlabel metal3 s 6882 40227 6980 40325 4 vdd
rlabel metal3 s 6882 39437 6980 39535 4 vdd
rlabel metal3 s 6882 41449 6980 41547 4 vdd
rlabel metal3 s 6450 38289 6548 38387 4 vdd
rlabel metal3 s 6882 43029 6980 43127 4 vdd
rlabel metal3 s 6882 40659 6980 40757 4 vdd
rlabel metal3 s 6450 43029 6548 43127 4 vdd
rlabel metal3 s 7660 40636 7758 40734 4 vdd
rlabel metal3 s 7660 43796 7758 43894 4 vdd
rlabel metal3 s 6450 39079 6548 39177 4 vdd
rlabel metal3 s 6882 42239 6980 42337 4 vdd
rlabel metal3 s 6450 42239 6548 42337 4 vdd
rlabel metal3 s 7660 40241 7758 40339 4 vdd
rlabel metal3 s 6450 37857 6548 37955 4 vdd
rlabel metal3 s 6882 38289 6980 38387 4 vdd
rlabel metal3 s 6882 39869 6980 39967 4 vdd
rlabel metal3 s 6882 43819 6980 43917 4 vdd
rlabel metal3 s 7660 43401 7758 43499 4 vdd
rlabel metal3 s 6450 41449 6548 41547 4 vdd
rlabel metal3 s 7660 41426 7758 41524 4 vdd
rlabel metal3 s 7660 42216 7758 42314 4 vdd
rlabel metal3 s 7660 39451 7758 39549 4 vdd
rlabel metal3 s 6882 43387 6980 43485 4 vdd
rlabel metal3 s 6450 43387 6548 43485 4 vdd
rlabel metal3 s 6450 38647 6548 38745 4 vdd
rlabel metal3 s 7264 38266 7362 38364 4 gnd
rlabel metal3 s 7264 43401 7362 43499 4 gnd
rlabel metal3 s 7264 40241 7362 40339 4 gnd
rlabel metal3 s 6450 41807 6548 41905 4 vdd
rlabel metal3 s 6450 41017 6548 41115 4 vdd
rlabel metal3 s 6450 40659 6548 40757 4 vdd
rlabel metal3 s 7660 41821 7758 41919 4 vdd
rlabel metal3 s 7264 42216 7362 42314 4 gnd
rlabel metal3 s 7264 39451 7362 39549 4 gnd
rlabel metal3 s 6450 42597 6548 42695 4 vdd
rlabel metal3 s 7660 39056 7758 39154 4 vdd
rlabel metal3 s 6882 39079 6980 39177 4 vdd
rlabel metal3 s 7264 40636 7362 40734 4 gnd
rlabel metal3 s 7264 41031 7362 41129 4 gnd
rlabel metal3 s 7264 43796 7362 43894 4 gnd
rlabel metal3 s 7264 39846 7362 39944 4 gnd
rlabel metal3 s 7264 37871 7362 37969 4 gnd
rlabel metal3 s 7264 42611 7362 42709 4 gnd
rlabel metal3 s 7264 39056 7362 39154 4 gnd
rlabel metal3 s 7264 41426 7362 41524 4 gnd
rlabel metal3 s 7264 43006 7362 43104 4 gnd
rlabel metal3 s 6882 41017 6980 41115 4 vdd
rlabel metal3 s 7264 38661 7362 38759 4 gnd
rlabel metal3 s 6882 38647 6980 38745 4 vdd
rlabel metal3 s 7264 41821 7362 41919 4 gnd
rlabel metal3 s 6882 42597 6980 42695 4 vdd
rlabel metal3 s 6882 37857 6980 37955 4 vdd
rlabel metal3 s 6450 39869 6548 39967 4 vdd
rlabel metal3 s 7660 38266 7758 38364 4 vdd
rlabel metal3 s 6025 39869 6123 39967 4 gnd
rlabel metal3 s 6025 41449 6123 41547 4 gnd
rlabel metal3 s 6025 47395 6123 47493 4 gnd
rlabel metal3 s 6025 50139 6123 50237 4 gnd
rlabel metal3 s 6025 47769 6123 47867 4 gnd
rlabel metal3 s 6025 42239 6123 42337 4 gnd
rlabel metal3 s 6025 45025 6123 45123 4 gnd
rlabel metal3 s 6025 48185 6123 48283 4 gnd
rlabel metal3 s 6025 38289 6123 38387 4 gnd
rlabel metal3 s 6025 42655 6123 42753 4 gnd
rlabel metal3 s 6025 44235 6123 44333 4 gnd
rlabel metal3 s 6025 39495 6123 39593 4 gnd
rlabel metal3 s 6025 44609 6123 44707 4 gnd
rlabel metal3 s 6025 40285 6123 40383 4 gnd
rlabel metal3 s 6025 43029 6123 43127 4 gnd
rlabel metal3 s 6025 43819 6123 43917 4 gnd
rlabel metal3 s 6025 48975 6123 49073 4 gnd
rlabel metal3 s 6025 38705 6123 38803 4 gnd
rlabel metal3 s 6025 46979 6123 47077 4 gnd
rlabel metal3 s 6025 43445 6123 43543 4 gnd
rlabel metal3 s 6025 45815 6123 45913 4 gnd
rlabel metal3 s 6025 37915 6123 38013 4 gnd
rlabel metal3 s 6025 40659 6123 40757 4 gnd
rlabel metal3 s 6025 41075 6123 41173 4 gnd
rlabel metal3 s 6025 48559 6123 48657 4 gnd
rlabel metal3 s 6025 41865 6123 41963 4 gnd
rlabel metal3 s 6025 45399 6123 45497 4 gnd
rlabel metal3 s 6025 39079 6123 39177 4 gnd
rlabel metal3 s 6025 49349 6123 49447 4 gnd
rlabel metal3 s 6025 49765 6123 49863 4 gnd
rlabel metal3 s 6025 46605 6123 46703 4 gnd
rlabel metal3 s 6025 46189 6123 46287 4 gnd
rlabel metal3 s 6025 29225 6123 29323 4 gnd
rlabel metal3 s 6025 32385 6123 32483 4 gnd
rlabel metal3 s 6025 35919 6123 36017 4 gnd
rlabel metal3 s 6025 31179 6123 31277 4 gnd
rlabel metal3 s 6025 26065 6123 26163 4 gnd
rlabel metal3 s 6025 28435 6123 28533 4 gnd
rlabel metal3 s 6025 32759 6123 32857 4 gnd
rlabel metal3 s 6025 28809 6123 28907 4 gnd
rlabel metal3 s 6025 33549 6123 33647 4 gnd
rlabel metal3 s 6025 30389 6123 30487 4 gnd
rlabel metal3 s 6025 31969 6123 32067 4 gnd
rlabel metal3 s 6025 27229 6123 27327 4 gnd
rlabel metal3 s 6025 33965 6123 34063 4 gnd
rlabel metal3 s 6025 36709 6123 36807 4 gnd
rlabel metal3 s 6025 25275 6123 25373 4 gnd
rlabel metal3 s 6025 27645 6123 27743 4 gnd
rlabel metal3 s 6025 37499 6123 37597 4 gnd
rlabel metal3 s 6025 25649 6123 25747 4 gnd
rlabel metal3 s 6025 26439 6123 26537 4 gnd
rlabel metal3 s 6025 35129 6123 35227 4 gnd
rlabel metal3 s 6025 37125 6123 37223 4 gnd
rlabel metal3 s 6025 29599 6123 29697 4 gnd
rlabel metal3 s 6025 30015 6123 30113 4 gnd
rlabel metal3 s 6025 35545 6123 35643 4 gnd
rlabel metal3 s 6025 30805 6123 30903 4 gnd
rlabel metal3 s 6025 34755 6123 34853 4 gnd
rlabel metal3 s 6025 34339 6123 34437 4 gnd
rlabel metal3 s 6025 36335 6123 36433 4 gnd
rlabel metal3 s 6025 31595 6123 31693 4 gnd
rlabel metal3 s 6025 28019 6123 28117 4 gnd
rlabel metal3 s 6025 33175 6123 33273 4 gnd
rlabel metal3 s 6025 26855 6123 26953 4 gnd
rlabel metal3 s 6450 35487 6548 35585 4 vdd
rlabel metal3 s 7264 36686 7362 36784 4 gnd
rlabel metal3 s 6882 32327 6980 32425 4 vdd
rlabel metal3 s 6450 36709 6548 36807 4 vdd
rlabel metal3 s 6882 36709 6980 36807 4 vdd
rlabel metal3 s 6450 33117 6548 33215 4 vdd
rlabel metal3 s 7660 37476 7758 37574 4 vdd
rlabel metal3 s 7264 32341 7362 32439 4 gnd
rlabel metal3 s 7264 37081 7362 37179 4 gnd
rlabel metal3 s 7660 31551 7758 31649 4 vdd
rlabel metal3 s 7264 35106 7362 35204 4 gnd
rlabel metal3 s 6882 31537 6980 31635 4 vdd
rlabel metal3 s 7660 31946 7758 32044 4 vdd
rlabel metal3 s 6450 33549 6548 33647 4 vdd
rlabel metal3 s 7660 35106 7758 35204 4 vdd
rlabel metal3 s 6450 36277 6548 36375 4 vdd
rlabel metal3 s 6450 31537 6548 31635 4 vdd
rlabel metal3 s 7264 37476 7362 37574 4 gnd
rlabel metal3 s 7660 32736 7758 32834 4 vdd
rlabel metal3 s 6882 35919 6980 36017 4 vdd
rlabel metal3 s 6450 37499 6548 37597 4 vdd
rlabel metal3 s 7264 34316 7362 34414 4 gnd
rlabel metal3 s 6882 34697 6980 34795 4 vdd
rlabel metal3 s 6882 35487 6980 35585 4 vdd
rlabel metal3 s 6450 32327 6548 32425 4 vdd
rlabel metal3 s 7660 33526 7758 33624 4 vdd
rlabel metal3 s 7264 31551 7362 31649 4 gnd
rlabel metal3 s 7660 32341 7758 32439 4 vdd
rlabel metal3 s 6450 34697 6548 34795 4 vdd
rlabel metal3 s 6450 32759 6548 32857 4 vdd
rlabel metal3 s 6882 31969 6980 32067 4 vdd
rlabel metal3 s 7660 37081 7758 37179 4 vdd
rlabel metal3 s 7264 35501 7362 35599 4 gnd
rlabel metal3 s 6882 33549 6980 33647 4 vdd
rlabel metal3 s 6450 33907 6548 34005 4 vdd
rlabel metal3 s 7660 33921 7758 34019 4 vdd
rlabel metal3 s 6882 33907 6980 34005 4 vdd
rlabel metal3 s 6450 35919 6548 36017 4 vdd
rlabel metal3 s 6882 37499 6980 37597 4 vdd
rlabel metal3 s 6882 37067 6980 37165 4 vdd
rlabel metal3 s 7660 33131 7758 33229 4 vdd
rlabel metal3 s 7660 34711 7758 34809 4 vdd
rlabel metal3 s 6450 34339 6548 34437 4 vdd
rlabel metal3 s 6882 33117 6980 33215 4 vdd
rlabel metal3 s 7660 36686 7758 36784 4 vdd
rlabel metal3 s 6882 32759 6980 32857 4 vdd
rlabel metal3 s 7264 31946 7362 32044 4 gnd
rlabel metal3 s 7264 35896 7362 35994 4 gnd
rlabel metal3 s 7660 34316 7758 34414 4 vdd
rlabel metal3 s 7264 33131 7362 33229 4 gnd
rlabel metal3 s 7264 33921 7362 34019 4 gnd
rlabel metal3 s 7660 35896 7758 35994 4 vdd
rlabel metal3 s 6450 37067 6548 37165 4 vdd
rlabel metal3 s 7660 35501 7758 35599 4 vdd
rlabel metal3 s 6882 36277 6980 36375 4 vdd
rlabel metal3 s 6450 31969 6548 32067 4 vdd
rlabel metal3 s 7264 36291 7362 36389 4 gnd
rlabel metal3 s 6450 35129 6548 35227 4 vdd
rlabel metal3 s 6882 35129 6980 35227 4 vdd
rlabel metal3 s 6882 34339 6980 34437 4 vdd
rlabel metal3 s 7660 36291 7758 36389 4 vdd
rlabel metal3 s 7264 34711 7362 34809 4 gnd
rlabel metal3 s 7264 33526 7362 33624 4 gnd
rlabel metal3 s 7264 32736 7362 32834 4 gnd
rlabel metal3 s 6882 25649 6980 25747 4 vdd
rlabel metal3 s 7660 31156 7758 31254 4 vdd
rlabel metal3 s 7660 30761 7758 30859 4 vdd
rlabel metal3 s 6882 28019 6980 28117 4 vdd
rlabel metal3 s 7660 26811 7758 26909 4 vdd
rlabel metal3 s 7660 28391 7758 28489 4 vdd
rlabel metal3 s 6450 30747 6548 30845 4 vdd
rlabel metal3 s 7264 26416 7362 26514 4 gnd
rlabel metal3 s 7264 27601 7362 27699 4 gnd
rlabel metal3 s 6450 30389 6548 30487 4 vdd
rlabel metal3 s 6450 31179 6548 31277 4 vdd
rlabel metal3 s 7264 26811 7362 26909 4 gnd
rlabel metal3 s 7660 25231 7758 25329 4 vdd
rlabel metal3 s 7660 29181 7758 29279 4 vdd
rlabel metal3 s 7264 25231 7362 25329 4 gnd
rlabel metal3 s 6882 28377 6980 28475 4 vdd
rlabel metal3 s 7264 29181 7362 29279 4 gnd
rlabel metal3 s 6882 28809 6980 28907 4 vdd
rlabel metal3 s 6450 26439 6548 26537 4 vdd
rlabel metal3 s 6882 27587 6980 27685 4 vdd
rlabel metal3 s 6450 27587 6548 27685 4 vdd
rlabel metal3 s 6450 25217 6548 25315 4 vdd
rlabel metal3 s 8092 25216 8190 25314 4 gnd
rlabel metal3 s 6450 27229 6548 27327 4 vdd
rlabel metal3 s 7660 27206 7758 27304 4 vdd
rlabel metal3 s 7264 26021 7362 26119 4 gnd
rlabel metal3 s 7264 30366 7362 30464 4 gnd
rlabel metal3 s 6450 25649 6548 25747 4 vdd
rlabel metal3 s 6882 29167 6980 29265 4 vdd
rlabel metal3 s 7264 29971 7362 30069 4 gnd
rlabel metal3 s 7264 27996 7362 28094 4 gnd
rlabel metal3 s 7264 31156 7362 31254 4 gnd
rlabel metal3 s 7660 29971 7758 30069 4 vdd
rlabel metal3 s 6450 28019 6548 28117 4 vdd
rlabel metal3 s 6882 26439 6980 26537 4 vdd
rlabel metal3 s 6882 25217 6980 25315 4 vdd
rlabel metal3 s 6450 26007 6548 26105 4 vdd
rlabel metal3 s 7660 26416 7758 26514 4 vdd
rlabel metal3 s 6450 26797 6548 26895 4 vdd
rlabel metal3 s 7264 27206 7362 27304 4 gnd
rlabel metal3 s 7660 25626 7758 25724 4 vdd
rlabel metal3 s 7660 27601 7758 27699 4 vdd
rlabel metal3 s 8517 25215 8615 25313 4 vdd
rlabel metal3 s 7660 27996 7758 28094 4 vdd
rlabel metal3 s 6450 29957 6548 30055 4 vdd
rlabel metal3 s 6450 29599 6548 29697 4 vdd
rlabel metal3 s 6882 27229 6980 27327 4 vdd
rlabel metal3 s 6450 29167 6548 29265 4 vdd
rlabel metal3 s 7264 28391 7362 28489 4 gnd
rlabel metal3 s 7660 29576 7758 29674 4 vdd
rlabel metal3 s 7660 30366 7758 30464 4 vdd
rlabel metal3 s 6882 31179 6980 31277 4 vdd
rlabel metal3 s 7660 28786 7758 28884 4 vdd
rlabel metal3 s 7264 28786 7362 28884 4 gnd
rlabel metal3 s 6450 28377 6548 28475 4 vdd
rlabel metal3 s 6882 26797 6980 26895 4 vdd
rlabel metal3 s 7264 30761 7362 30859 4 gnd
rlabel metal3 s 6882 30389 6980 30487 4 vdd
rlabel metal3 s 7660 26021 7758 26119 4 vdd
rlabel metal3 s 7264 29576 7362 29674 4 gnd
rlabel metal3 s 6882 26007 6980 26105 4 vdd
rlabel metal3 s 6450 28809 6548 28907 4 vdd
rlabel metal3 s 6882 29599 6980 29697 4 vdd
rlabel metal3 s 6882 30747 6980 30845 4 vdd
rlabel metal3 s 6882 29957 6980 30055 4 vdd
rlabel metal3 s 7264 25626 7362 25724 4 gnd
rlabel metal3 s 9560 25231 9658 25329 4 gnd
rlabel metal3 s 11208 25231 11306 25329 4 vdd
rlabel metal3 s 1156 5086 1254 5184 4 gnd
rlabel metal3 s 7660 24441 7758 24539 4 vdd
rlabel metal3 s 6450 24069 6548 24167 4 vdd
rlabel metal3 s 7660 24836 7758 24934 4 vdd
rlabel metal3 s 6450 19687 6548 19785 4 vdd
rlabel metal3 s 6882 21699 6980 21797 4 vdd
rlabel metal3 s 6882 24859 6980 24957 4 vdd
rlabel metal3 s 7660 20096 7758 20194 4 vdd
rlabel metal3 s 6450 21267 6548 21365 4 vdd
rlabel metal3 s 6882 18897 6980 18995 4 vdd
rlabel metal3 s 7660 18911 7758 19009 4 vdd
rlabel metal3 s 6882 20909 6980 21007 4 vdd
rlabel metal3 s 6450 20909 6548 21007 4 vdd
rlabel metal3 s 6882 20477 6980 20575 4 vdd
rlabel metal3 s 6882 24069 6980 24167 4 vdd
rlabel metal3 s 7660 22071 7758 22169 4 vdd
rlabel metal3 s 7660 23256 7758 23354 4 vdd
rlabel metal3 s 6450 20119 6548 20217 4 vdd
rlabel metal3 s 7264 20096 7362 20194 4 gnd
rlabel metal3 s 7264 24046 7362 24144 4 gnd
rlabel metal3 s 6882 22847 6980 22945 4 vdd
rlabel metal3 s 7660 19306 7758 19404 4 vdd
rlabel metal3 s 6450 23279 6548 23377 4 vdd
rlabel metal3 s 7264 23651 7362 23749 4 gnd
rlabel metal3 s 7660 22861 7758 22959 4 vdd
rlabel metal3 s 7660 20491 7758 20589 4 vdd
rlabel metal3 s 7264 19306 7362 19404 4 gnd
rlabel metal3 s 7264 21676 7362 21774 4 gnd
rlabel metal3 s 7264 22071 7362 22169 4 gnd
rlabel metal3 s 7264 20491 7362 20589 4 gnd
rlabel metal3 s 6450 24427 6548 24525 4 vdd
rlabel metal3 s 7264 24441 7362 24539 4 gnd
rlabel metal3 s 7264 22861 7362 22959 4 gnd
rlabel metal3 s 6450 22489 6548 22587 4 vdd
rlabel metal3 s 6450 20477 6548 20575 4 vdd
rlabel metal3 s 7660 24046 7758 24144 4 vdd
rlabel metal3 s 7660 21281 7758 21379 4 vdd
rlabel metal3 s 7264 24836 7362 24934 4 gnd
rlabel metal3 s 7264 23256 7362 23354 4 gnd
rlabel metal3 s 7660 20886 7758 20984 4 vdd
rlabel metal3 s 6450 22057 6548 22155 4 vdd
rlabel metal3 s 7264 21281 7362 21379 4 gnd
rlabel metal3 s 7660 23651 7758 23749 4 vdd
rlabel metal3 s 6450 21699 6548 21797 4 vdd
rlabel metal3 s 6882 24427 6980 24525 4 vdd
rlabel metal3 s 7660 19701 7758 19799 4 vdd
rlabel metal3 s 7660 22466 7758 22564 4 vdd
rlabel metal3 s 6450 24859 6548 24957 4 vdd
rlabel metal3 s 6882 23279 6980 23377 4 vdd
rlabel metal3 s 6882 22489 6980 22587 4 vdd
rlabel metal3 s 7264 22466 7362 22564 4 gnd
rlabel metal3 s 7264 19701 7362 19799 4 gnd
rlabel metal3 s 6450 18897 6548 18995 4 vdd
rlabel metal3 s 6882 19687 6980 19785 4 vdd
rlabel metal3 s 6450 19329 6548 19427 4 vdd
rlabel metal3 s 6450 22847 6548 22945 4 vdd
rlabel metal3 s 7264 20886 7362 20984 4 gnd
rlabel metal3 s 6882 22057 6980 22155 4 vdd
rlabel metal3 s 6882 19329 6980 19427 4 vdd
rlabel metal3 s 6882 20119 6980 20217 4 vdd
rlabel metal3 s 7264 18911 7362 19009 4 gnd
rlabel metal3 s 6450 23637 6548 23735 4 vdd
rlabel metal3 s 6882 23637 6980 23735 4 vdd
rlabel metal3 s 7660 21676 7758 21774 4 vdd
rlabel metal3 s 6882 21267 6980 21365 4 vdd
rlabel metal3 s 7264 18516 7362 18614 4 gnd
rlabel metal3 s 6450 14157 6548 14255 4 vdd
rlabel metal3 s 7660 17726 7758 17824 4 vdd
rlabel metal3 s 7264 17726 7362 17824 4 gnd
rlabel metal3 s 7264 15751 7362 15849 4 gnd
rlabel metal3 s 7264 14566 7362 14664 4 gnd
rlabel metal3 s 7264 16936 7362 17034 4 gnd
rlabel metal3 s 6882 17749 6980 17847 4 vdd
rlabel metal3 s 6882 18539 6980 18637 4 vdd
rlabel metal3 s 6882 12577 6980 12675 4 vdd
rlabel metal3 s 6450 17317 6548 17415 4 vdd
rlabel metal3 s 6882 14947 6980 15045 4 vdd
rlabel metal3 s 6450 17749 6548 17847 4 vdd
rlabel metal3 s 7660 15356 7758 15454 4 vdd
rlabel metal3 s 6450 13799 6548 13897 4 vdd
rlabel metal3 s 6450 13367 6548 13465 4 vdd
rlabel metal3 s 6450 16169 6548 16267 4 vdd
rlabel metal3 s 6882 14589 6980 14687 4 vdd
rlabel metal3 s 7660 18516 7758 18614 4 vdd
rlabel metal3 s 7660 14171 7758 14269 4 vdd
rlabel metal3 s 7264 15356 7362 15454 4 gnd
rlabel metal3 s 6450 14589 6548 14687 4 vdd
rlabel metal3 s 6450 13009 6548 13107 4 vdd
rlabel metal3 s 7264 13776 7362 13874 4 gnd
rlabel metal3 s 6450 14947 6548 15045 4 vdd
rlabel metal3 s 7264 14961 7362 15059 4 gnd
rlabel metal3 s 7660 14961 7758 15059 4 vdd
rlabel metal3 s 7660 16936 7758 17034 4 vdd
rlabel metal3 s 6450 18107 6548 18205 4 vdd
rlabel metal3 s 6882 13009 6980 13107 4 vdd
rlabel metal3 s 6882 13367 6980 13465 4 vdd
rlabel metal3 s 7264 17331 7362 17429 4 gnd
rlabel metal3 s 6882 15737 6980 15835 4 vdd
rlabel metal3 s 6882 13799 6980 13897 4 vdd
rlabel metal3 s 6450 12577 6548 12675 4 vdd
rlabel metal3 s 7660 12986 7758 13084 4 vdd
rlabel metal3 s 6882 15379 6980 15477 4 vdd
rlabel metal3 s 7660 16146 7758 16244 4 vdd
rlabel metal3 s 7660 18121 7758 18219 4 vdd
rlabel metal3 s 7660 12591 7758 12689 4 vdd
rlabel metal3 s 7660 14566 7758 14664 4 vdd
rlabel metal3 s 6882 16169 6980 16267 4 vdd
rlabel metal3 s 7264 16146 7362 16244 4 gnd
rlabel metal3 s 7264 13381 7362 13479 4 gnd
rlabel metal3 s 6450 16527 6548 16625 4 vdd
rlabel metal3 s 7660 17331 7758 17429 4 vdd
rlabel metal3 s 6882 18107 6980 18205 4 vdd
rlabel metal3 s 6882 16959 6980 17057 4 vdd
rlabel metal3 s 7264 12986 7362 13084 4 gnd
rlabel metal3 s 7660 13776 7758 13874 4 vdd
rlabel metal3 s 7264 16541 7362 16639 4 gnd
rlabel metal3 s 6450 16959 6548 17057 4 vdd
rlabel metal3 s 6450 15379 6548 15477 4 vdd
rlabel metal3 s 7264 14171 7362 14269 4 gnd
rlabel metal3 s 7660 16541 7758 16639 4 vdd
rlabel metal3 s 6450 18539 6548 18637 4 vdd
rlabel metal3 s 6882 16527 6980 16625 4 vdd
rlabel metal3 s 6882 17317 6980 17415 4 vdd
rlabel metal3 s 6450 15737 6548 15835 4 vdd
rlabel metal3 s 7264 18121 7362 18219 4 gnd
rlabel metal3 s 7660 15751 7758 15849 4 vdd
rlabel metal3 s 7264 12591 7362 12689 4 gnd
rlabel metal3 s 6882 14157 6980 14255 4 vdd
rlabel metal3 s 7660 13381 7758 13479 4 vdd
rlabel metal3 s 6025 15379 6123 15477 4 gnd
rlabel metal3 s 6025 21699 6123 21797 4 gnd
rlabel metal3 s 6025 16169 6123 16267 4 gnd
rlabel metal3 s 6025 24069 6123 24167 4 gnd
rlabel metal3 s 6025 13425 6123 13523 4 gnd
rlabel metal3 s 6025 23279 6123 23377 4 gnd
rlabel metal3 s 6025 24485 6123 24583 4 gnd
rlabel metal3 s 6025 15795 6123 15893 4 gnd
rlabel metal3 s 6025 19745 6123 19843 4 gnd
rlabel metal3 s 6025 17375 6123 17473 4 gnd
rlabel metal3 s 6025 16959 6123 17057 4 gnd
rlabel metal3 s 6025 15005 6123 15103 4 gnd
rlabel metal3 s 6025 20535 6123 20633 4 gnd
rlabel metal3 s 6025 22905 6123 23003 4 gnd
rlabel metal3 s 6025 14589 6123 14687 4 gnd
rlabel metal3 s 6025 22489 6123 22587 4 gnd
rlabel metal3 s 6025 21325 6123 21423 4 gnd
rlabel metal3 s 6025 24859 6123 24957 4 gnd
rlabel metal3 s 6025 17749 6123 17847 4 gnd
rlabel metal3 s 6025 12635 6123 12733 4 gnd
rlabel metal3 s 6025 19329 6123 19427 4 gnd
rlabel metal3 s 6025 20909 6123 21007 4 gnd
rlabel metal3 s 6025 16585 6123 16683 4 gnd
rlabel metal3 s 6025 23695 6123 23793 4 gnd
rlabel metal3 s 6025 13799 6123 13897 4 gnd
rlabel metal3 s 6025 13009 6123 13107 4 gnd
rlabel metal3 s 6025 14215 6123 14313 4 gnd
rlabel metal3 s 6025 18539 6123 18637 4 gnd
rlabel metal3 s 6025 20119 6123 20217 4 gnd
rlabel metal3 s 6025 18955 6123 19053 4 gnd
rlabel metal3 s 6025 22115 6123 22213 4 gnd
rlabel metal3 s 6025 18165 6123 18263 4 gnd
rlabel metal3 s 6025 3945 6123 4043 4 gnd
rlabel metal3 s 3046 3513 3144 3611 4 gnd
rlabel metal3 s 3850 1136 3948 1234 4 gnd
rlabel metal3 s 4246 1136 4344 1234 4 vdd
rlabel metal3 s 6025 1575 6123 1673 4 gnd
rlabel metal3 s 6025 11845 6123 11943 4 gnd
rlabel metal3 s 2611 7479 2709 7577 4 gnd
rlabel metal3 s 3036 6689 3134 6787 4 vdd
rlabel metal3 s 1752 346 1850 444 4 gnd
rlabel metal3 s 2148 2716 2246 2814 4 vdd
rlabel metal3 s 6025 3155 6123 3253 4 gnd
rlabel metal3 s 3471 1143 3569 1241 4 vdd
rlabel metal3 s 3468 7479 3566 7577 4 vdd
rlabel metal3 s 3850 6666 3948 6764 4 gnd
rlabel metal3 s 6025 5109 6123 5207 4 gnd
rlabel metal3 s 6025 12219 6123 12317 4 gnd
rlabel metal3 s 6025 11055 6123 11153 4 gnd
rlabel metal3 s 6025 369 6123 467 4 gnd
rlabel metal3 s 6025 6315 6123 6413 4 gnd
rlabel metal3 s 4246 6666 4344 6764 4 vdd
rlabel metal3 s 3468 6689 3566 6787 4 vdd
rlabel metal3 s 2148 346 2246 444 4 vdd
rlabel metal3 s 1752 2716 1850 2814 4 gnd
rlabel metal3 s 4246 2716 4344 2814 4 vdd
rlabel metal3 s 6025 10265 6123 10363 4 gnd
rlabel metal3 s 6025 10639 6123 10737 4 gnd
rlabel metal3 s 4246 5086 4344 5184 4 vdd
rlabel metal3 s 6025 9475 6123 9573 4 gnd
rlabel metal3 s 3850 7456 3948 7554 4 gnd
rlabel metal3 s 3046 2723 3144 2821 4 gnd
rlabel metal3 s 6025 1949 6123 2047 4 gnd
rlabel metal3 s 6025 2365 6123 2463 4 gnd
rlabel metal3 s 3850 5876 3948 5974 4 gnd
rlabel metal3 s 3036 5109 3134 5207 4 vdd
rlabel metal3 s 4246 346 4344 444 4 vdd
rlabel metal3 s 6025 4319 6123 4417 4 gnd
rlabel metal3 s 1552 5086 1650 5184 4 vdd
rlabel metal3 s 6025 4735 6123 4833 4 gnd
rlabel metal3 s 3046 1143 3144 1241 4 gnd
rlabel metal3 s 3471 353 3569 451 4 vdd
rlabel metal3 s 6025 7479 6123 7577 4 gnd
rlabel metal3 s 6025 11429 6123 11527 4 gnd
rlabel metal3 s 6025 785 6123 883 4 gnd
rlabel metal3 s 6025 9059 6123 9157 4 gnd
rlabel metal3 s 3046 353 3144 451 4 gnd
rlabel metal3 s 6025 9849 6123 9947 4 gnd
rlabel metal3 s 3036 5899 3134 5997 4 vdd
rlabel metal3 s 6025 8269 6123 8367 4 gnd
rlabel metal3 s 3036 7479 3134 7577 4 vdd
rlabel metal3 s 3471 3513 3569 3611 4 vdd
rlabel metal3 s 6025 5899 6123 5997 4 gnd
rlabel metal3 s 6025 7105 6123 7203 4 gnd
rlabel metal3 s 2611 6689 2709 6787 4 gnd
rlabel metal3 s 6025 6689 6123 6787 4 gnd
rlabel metal3 s 3468 5899 3566 5997 4 vdd
rlabel metal3 s 3850 346 3948 444 4 gnd
rlabel metal3 s 6025 1159 6123 1257 4 gnd
rlabel metal3 s 2611 5899 2709 5997 4 gnd
rlabel metal3 s 4246 3506 4344 3604 4 vdd
rlabel metal3 s 4246 7456 4344 7554 4 vdd
rlabel metal3 s 3468 5109 3566 5207 4 vdd
rlabel metal3 s 6025 3529 6123 3627 4 gnd
rlabel metal3 s 3471 2723 3569 2821 4 vdd
rlabel metal3 s 4246 5876 4344 5974 4 vdd
rlabel metal3 s 6025 7895 6123 7993 4 gnd
rlabel metal3 s 2611 5109 2709 5207 4 gnd
rlabel metal3 s 3850 3506 3948 3604 4 gnd
rlabel metal3 s 6025 5525 6123 5623 4 gnd
rlabel metal3 s 3850 5086 3948 5184 4 gnd
rlabel metal3 s 3850 2716 3948 2814 4 gnd
rlabel metal3 s 6025 8685 6123 8783 4 gnd
rlabel metal3 s 6025 2739 6123 2837 4 gnd
rlabel metal3 s 7660 12196 7758 12294 4 vdd
rlabel metal3 s 6882 11429 6980 11527 4 vdd
rlabel metal3 s 6882 7047 6980 7145 4 vdd
rlabel metal3 s 7264 9431 7362 9529 4 gnd
rlabel metal3 s 7264 9036 7362 9134 4 gnd
rlabel metal3 s 6450 9849 6548 9947 4 vdd
rlabel metal3 s 6882 6689 6980 6787 4 vdd
rlabel metal3 s 7660 8246 7758 8344 4 vdd
rlabel metal3 s 7264 10221 7362 10319 4 gnd
rlabel metal3 s 6882 7837 6980 7935 4 vdd
rlabel metal3 s 7264 7456 7362 7554 4 gnd
rlabel metal3 s 7264 6666 7362 6764 4 gnd
rlabel metal3 s 6882 8269 6980 8367 4 vdd
rlabel metal3 s 6882 9417 6980 9515 4 vdd
rlabel metal3 s 7660 7456 7758 7554 4 vdd
rlabel metal3 s 7660 9036 7758 9134 4 vdd
rlabel metal3 s 6882 9849 6980 9947 4 vdd
rlabel metal3 s 6450 7479 6548 7577 4 vdd
rlabel metal3 s 6450 8269 6548 8367 4 vdd
rlabel metal3 s 7660 8641 7758 8739 4 vdd
rlabel metal3 s 6450 10997 6548 11095 4 vdd
rlabel metal3 s 6450 6689 6548 6787 4 vdd
rlabel metal3 s 6450 12219 6548 12317 4 vdd
rlabel metal3 s 6450 9059 6548 9157 4 vdd
rlabel metal3 s 7660 9826 7758 9924 4 vdd
rlabel metal3 s 6450 7837 6548 7935 4 vdd
rlabel metal3 s 7660 11801 7758 11899 4 vdd
rlabel metal3 s 7660 11011 7758 11109 4 vdd
rlabel metal3 s 6882 7479 6980 7577 4 vdd
rlabel metal3 s 7660 11406 7758 11504 4 vdd
rlabel metal3 s 7660 9431 7758 9529 4 vdd
rlabel metal3 s 6450 11787 6548 11885 4 vdd
rlabel metal3 s 7264 11011 7362 11109 4 gnd
rlabel metal3 s 6882 6257 6980 6355 4 vdd
rlabel metal3 s 6450 11429 6548 11527 4 vdd
rlabel metal3 s 7660 6666 7758 6764 4 vdd
rlabel metal3 s 7660 7851 7758 7949 4 vdd
rlabel metal3 s 6450 7047 6548 7145 4 vdd
rlabel metal3 s 7264 7851 7362 7949 4 gnd
rlabel metal3 s 7264 10616 7362 10714 4 gnd
rlabel metal3 s 6882 12219 6980 12317 4 vdd
rlabel metal3 s 6882 10207 6980 10305 4 vdd
rlabel metal3 s 7264 8641 7362 8739 4 gnd
rlabel metal3 s 6450 8627 6548 8725 4 vdd
rlabel metal3 s 6450 10639 6548 10737 4 vdd
rlabel metal3 s 7264 9826 7362 9924 4 gnd
rlabel metal3 s 6882 10997 6980 11095 4 vdd
rlabel metal3 s 7660 10616 7758 10714 4 vdd
rlabel metal3 s 7264 11801 7362 11899 4 gnd
rlabel metal3 s 7264 8246 7362 8344 4 gnd
rlabel metal3 s 6882 8627 6980 8725 4 vdd
rlabel metal3 s 6450 10207 6548 10305 4 vdd
rlabel metal3 s 7660 7061 7758 7159 4 vdd
rlabel metal3 s 6450 9417 6548 9515 4 vdd
rlabel metal3 s 7660 6271 7758 6369 4 vdd
rlabel metal3 s 6882 10639 6980 10737 4 vdd
rlabel metal3 s 6882 11787 6980 11885 4 vdd
rlabel metal3 s 7264 7061 7362 7159 4 gnd
rlabel metal3 s 7660 10221 7758 10319 4 vdd
rlabel metal3 s 7264 12196 7362 12294 4 gnd
rlabel metal3 s 7264 6271 7362 6369 4 gnd
rlabel metal3 s 7264 11406 7362 11504 4 gnd
rlabel metal3 s 6882 9059 6980 9157 4 vdd
rlabel metal3 s 6450 6257 6548 6355 4 vdd
rlabel metal3 s 6450 4677 6548 4775 4 vdd
rlabel metal3 s 6450 5109 6548 5207 4 vdd
rlabel metal3 s 7660 3111 7758 3209 4 vdd
rlabel metal3 s 7660 3901 7758 3999 4 vdd
rlabel metal3 s 6450 4319 6548 4417 4 vdd
rlabel metal3 s 7264 4296 7362 4394 4 gnd
rlabel metal3 s 7660 5481 7758 5579 4 vdd
rlabel metal3 s 6450 727 6548 825 4 vdd
rlabel metal3 s 6882 1159 6980 1257 4 vdd
rlabel metal3 s 6450 369 6548 467 4 vdd
rlabel metal3 s 6882 2739 6980 2837 4 vdd
rlabel metal3 s 7660 741 7758 839 4 vdd
rlabel metal3 s 7264 3901 7362 3999 4 gnd
rlabel metal3 s 6450 5467 6548 5565 4 vdd
rlabel metal3 s 7264 3111 7362 3209 4 gnd
rlabel metal3 s 7264 741 7362 839 4 gnd
rlabel metal3 s 7660 3506 7758 3604 4 vdd
rlabel metal3 s 6882 1517 6980 1615 4 vdd
rlabel metal3 s 7264 1136 7362 1234 4 gnd
rlabel metal3 s 6450 1949 6548 2047 4 vdd
rlabel metal3 s 7264 3506 7362 3604 4 gnd
rlabel metal3 s 6882 5467 6980 5565 4 vdd
rlabel metal3 s 7660 5876 7758 5974 4 vdd
rlabel metal3 s 6882 4677 6980 4775 4 vdd
rlabel metal3 s 7660 2716 7758 2814 4 vdd
rlabel metal3 s 7264 1531 7362 1629 4 gnd
rlabel metal3 s 7660 5086 7758 5184 4 vdd
rlabel metal3 s 6882 3097 6980 3195 4 vdd
rlabel metal3 s 6450 3097 6548 3195 4 vdd
rlabel metal3 s 7264 1926 7362 2024 4 gnd
rlabel metal3 s 6882 3887 6980 3985 4 vdd
rlabel metal3 s 6882 2307 6980 2405 4 vdd
rlabel metal3 s 6450 3887 6548 3985 4 vdd
rlabel metal3 s 6450 1159 6548 1257 4 vdd
rlabel metal3 s 7660 4296 7758 4394 4 vdd
rlabel metal3 s 8517 -234 8615 -136 4 vdd
rlabel metal3 s 6882 369 6980 467 4 vdd
rlabel metal3 s 7660 1136 7758 1234 4 vdd
rlabel metal3 s 7685 -240 7783 -142 4 vdd
rlabel metal3 s 7264 5481 7362 5579 4 gnd
rlabel metal3 s 7660 346 7758 444 4 vdd
rlabel metal3 s 7660 4691 7758 4789 4 vdd
rlabel metal3 s 6450 2307 6548 2405 4 vdd
rlabel metal3 s 7264 346 7362 444 4 gnd
rlabel metal3 s 6450 2739 6548 2837 4 vdd
rlabel metal3 s 6882 727 6980 825 4 vdd
rlabel metal3 s 7264 4691 7362 4789 4 gnd
rlabel metal3 s 7264 2321 7362 2419 4 gnd
rlabel metal3 s 6450 1517 6548 1615 4 vdd
rlabel metal3 s 6882 1949 6980 2047 4 vdd
rlabel metal3 s 6450 5899 6548 5997 4 vdd
rlabel metal3 s 7660 1926 7758 2024 4 vdd
rlabel metal3 s 6882 4319 6980 4417 4 vdd
rlabel metal3 s 7660 2321 7758 2419 4 vdd
rlabel metal3 s 7660 1531 7758 1629 4 vdd
rlabel metal3 s 7264 2716 7362 2814 4 gnd
rlabel metal3 s 7264 5086 7362 5184 4 gnd
rlabel metal3 s 6450 3529 6548 3627 4 vdd
rlabel metal3 s 6882 3529 6980 3627 4 vdd
rlabel metal3 s 6882 5899 6980 5997 4 vdd
rlabel metal3 s 7264 5876 7362 5974 4 gnd
rlabel metal3 s 6882 5109 6980 5207 4 vdd
rlabel metal3 s 11208 -246 11306 -148 4 vdd
rlabel metal2 s 7960 -313 7988 -285 4 wl_en
rlabel metal1 s 19 0 47 7900 4 addr_0
rlabel metal1 s 99 0 127 7900 4 addr_1
rlabel metal1 s 179 0 207 7900 4 addr_2
rlabel metal1 s 259 0 287 7900 4 addr_3
rlabel metal1 s 339 0 367 7900 4 addr_4
rlabel metal1 s 419 0 447 7900 4 addr_5
rlabel metal1 s 499 0 527 7900 4 addr_6
rlabel locali s 11979 25400 11979 25400 4 wl_64
rlabel locali s 11979 25950 11979 25950 4 wl_65
rlabel locali s 11979 26190 11979 26190 4 wl_66
rlabel locali s 11979 26740 11979 26740 4 wl_67
rlabel locali s 11979 26980 11979 26980 4 wl_68
rlabel locali s 11979 27530 11979 27530 4 wl_69
rlabel locali s 11979 27770 11979 27770 4 wl_70
rlabel locali s 11979 28320 11979 28320 4 wl_71
rlabel locali s 11979 28560 11979 28560 4 wl_72
rlabel locali s 11979 29110 11979 29110 4 wl_73
rlabel locali s 11979 29350 11979 29350 4 wl_74
rlabel locali s 11979 29900 11979 29900 4 wl_75
rlabel locali s 11979 30140 11979 30140 4 wl_76
rlabel locali s 11979 30690 11979 30690 4 wl_77
rlabel locali s 11979 30930 11979 30930 4 wl_78
rlabel locali s 11979 31480 11979 31480 4 wl_79
rlabel locali s 11979 31720 11979 31720 4 wl_80
rlabel locali s 11979 32270 11979 32270 4 wl_81
rlabel locali s 11979 32510 11979 32510 4 wl_82
rlabel locali s 11979 33060 11979 33060 4 wl_83
rlabel locali s 11979 33300 11979 33300 4 wl_84
rlabel locali s 11979 33850 11979 33850 4 wl_85
rlabel locali s 11979 34090 11979 34090 4 wl_86
rlabel locali s 11979 34640 11979 34640 4 wl_87
rlabel locali s 11979 34880 11979 34880 4 wl_88
rlabel locali s 11979 35430 11979 35430 4 wl_89
rlabel locali s 11979 35670 11979 35670 4 wl_90
rlabel locali s 11979 36220 11979 36220 4 wl_91
rlabel locali s 11979 36460 11979 36460 4 wl_92
rlabel locali s 11979 37010 11979 37010 4 wl_93
rlabel locali s 11979 37250 11979 37250 4 wl_94
rlabel locali s 11979 37800 11979 37800 4 wl_95
rlabel locali s 11979 38040 11979 38040 4 wl_96
rlabel locali s 11979 38590 11979 38590 4 wl_97
rlabel locali s 11979 38830 11979 38830 4 wl_98
rlabel locali s 11979 39380 11979 39380 4 wl_99
rlabel locali s 11979 39620 11979 39620 4 wl_100
rlabel locali s 11979 40170 11979 40170 4 wl_101
rlabel locali s 11979 40410 11979 40410 4 wl_102
rlabel locali s 11979 40960 11979 40960 4 wl_103
rlabel locali s 11979 41200 11979 41200 4 wl_104
rlabel locali s 11979 41750 11979 41750 4 wl_105
rlabel locali s 11979 41990 11979 41990 4 wl_106
rlabel locali s 11979 42540 11979 42540 4 wl_107
rlabel locali s 11979 42780 11979 42780 4 wl_108
rlabel locali s 11979 43330 11979 43330 4 wl_109
rlabel locali s 11979 43570 11979 43570 4 wl_110
rlabel locali s 11979 44120 11979 44120 4 wl_111
rlabel locali s 11979 44360 11979 44360 4 wl_112
rlabel locali s 11979 44910 11979 44910 4 wl_113
rlabel locali s 11979 45150 11979 45150 4 wl_114
rlabel locali s 11979 45700 11979 45700 4 wl_115
rlabel locali s 11979 45940 11979 45940 4 wl_116
rlabel locali s 11979 46490 11979 46490 4 wl_117
rlabel locali s 11979 46730 11979 46730 4 wl_118
rlabel locali s 11979 47280 11979 47280 4 wl_119
rlabel locali s 11979 47520 11979 47520 4 wl_120
rlabel locali s 11979 48070 11979 48070 4 wl_121
rlabel locali s 11979 48310 11979 48310 4 wl_122
rlabel locali s 11979 48860 11979 48860 4 wl_123
rlabel locali s 11979 49100 11979 49100 4 wl_124
rlabel locali s 11979 49650 11979 49650 4 wl_125
rlabel locali s 11979 49890 11979 49890 4 wl_126
rlabel locali s 11979 50440 11979 50440 4 wl_127
rlabel locali s 10784 -120 10784 -120 4 rbl_wl
rlabel locali s 11979 670 11979 670 4 wl_1
rlabel locali s 11979 910 11979 910 4 wl_2
rlabel locali s 11979 1460 11979 1460 4 wl_3
rlabel locali s 11979 1700 11979 1700 4 wl_4
rlabel locali s 11979 2250 11979 2250 4 wl_5
rlabel locali s 11979 2490 11979 2490 4 wl_6
rlabel locali s 11979 3040 11979 3040 4 wl_7
rlabel locali s 11979 3280 11979 3280 4 wl_8
rlabel locali s 11979 3830 11979 3830 4 wl_9
rlabel locali s 11979 4070 11979 4070 4 wl_10
rlabel locali s 11979 4620 11979 4620 4 wl_11
rlabel locali s 11979 4860 11979 4860 4 wl_12
rlabel locali s 11979 5410 11979 5410 4 wl_13
rlabel locali s 11979 5650 11979 5650 4 wl_14
rlabel locali s 11979 6200 11979 6200 4 wl_15
rlabel locali s 11979 6440 11979 6440 4 wl_16
rlabel locali s 11979 6990 11979 6990 4 wl_17
rlabel locali s 11979 7230 11979 7230 4 wl_18
rlabel locali s 11979 7780 11979 7780 4 wl_19
rlabel locali s 11979 8020 11979 8020 4 wl_20
rlabel locali s 11979 8570 11979 8570 4 wl_21
rlabel locali s 11979 8810 11979 8810 4 wl_22
rlabel locali s 11979 9360 11979 9360 4 wl_23
rlabel locali s 11979 9600 11979 9600 4 wl_24
rlabel locali s 11979 10150 11979 10150 4 wl_25
rlabel locali s 11979 10390 11979 10390 4 wl_26
rlabel locali s 11979 10940 11979 10940 4 wl_27
rlabel locali s 11979 11180 11979 11180 4 wl_28
rlabel locali s 11979 11730 11979 11730 4 wl_29
rlabel locali s 11979 11970 11979 11970 4 wl_30
rlabel locali s 11979 12520 11979 12520 4 wl_31
rlabel locali s 11979 12760 11979 12760 4 wl_32
rlabel locali s 11979 13310 11979 13310 4 wl_33
rlabel locali s 11979 13550 11979 13550 4 wl_34
rlabel locali s 11979 14100 11979 14100 4 wl_35
rlabel locali s 11979 14340 11979 14340 4 wl_36
rlabel locali s 11979 14890 11979 14890 4 wl_37
rlabel locali s 11979 15130 11979 15130 4 wl_38
rlabel locali s 11979 15680 11979 15680 4 wl_39
rlabel locali s 11979 15920 11979 15920 4 wl_40
rlabel locali s 11979 16470 11979 16470 4 wl_41
rlabel locali s 11979 16710 11979 16710 4 wl_42
rlabel locali s 11979 17260 11979 17260 4 wl_43
rlabel locali s 11979 17500 11979 17500 4 wl_44
rlabel locali s 11979 18050 11979 18050 4 wl_45
rlabel locali s 11979 18290 11979 18290 4 wl_46
rlabel locali s 11979 18840 11979 18840 4 wl_47
rlabel locali s 11979 19080 11979 19080 4 wl_48
rlabel locali s 11979 19630 11979 19630 4 wl_49
rlabel locali s 11979 19870 11979 19870 4 wl_50
rlabel locali s 11979 20420 11979 20420 4 wl_51
rlabel locali s 11979 20660 11979 20660 4 wl_52
rlabel locali s 11979 21210 11979 21210 4 wl_53
rlabel locali s 11979 21450 11979 21450 4 wl_54
rlabel locali s 11979 22000 11979 22000 4 wl_55
rlabel locali s 11979 22240 11979 22240 4 wl_56
rlabel locali s 11979 22790 11979 22790 4 wl_57
rlabel locali s 11979 23030 11979 23030 4 wl_58
rlabel locali s 11979 23580 11979 23580 4 wl_59
rlabel locali s 11979 23820 11979 23820 4 wl_60
rlabel locali s 11979 24370 11979 24370 4 wl_61
rlabel locali s 11979 24610 11979 24610 4 wl_62
rlabel locali s 11979 25160 11979 25160 4 wl_63
rlabel locali s 11979 120 11979 120 4 wl_0
<< properties >>
string FIXED_BBOX 7945 -332 8003 -331
string GDS_END 6670770
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 6475980
<< end >>
