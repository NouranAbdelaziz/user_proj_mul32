magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< locali >>
rect 1181 8861 1215 8877
rect 1181 8811 1215 8827
rect 11165 8861 11199 8877
rect 11165 8811 11199 8827
rect 21149 8861 21183 8877
rect 21149 8811 21183 8827
rect 31133 8861 31167 8877
rect 31133 8811 31167 8827
<< viali >>
rect 1181 8827 1215 8861
rect 11165 8827 11199 8861
rect 21149 8827 21183 8861
rect 31133 8827 31167 8861
<< metal1 >>
rect 1169 8861 1227 8867
rect 1169 8827 1181 8861
rect 1215 8858 1227 8861
rect 9967 8858 9973 8870
rect 1215 8830 9973 8858
rect 1215 8827 1227 8830
rect 1169 8821 1227 8827
rect 9967 8818 9973 8830
rect 10025 8818 10031 8870
rect 11153 8861 11211 8867
rect 11153 8827 11165 8861
rect 11199 8858 11211 8861
rect 19951 8858 19957 8870
rect 11199 8830 19957 8858
rect 11199 8827 11211 8830
rect 11153 8821 11211 8827
rect 19951 8818 19957 8830
rect 20009 8818 20015 8870
rect 21137 8861 21195 8867
rect 21137 8827 21149 8861
rect 21183 8858 21195 8861
rect 29935 8858 29941 8870
rect 21183 8830 29941 8858
rect 21183 8827 21195 8830
rect 21137 8821 21195 8827
rect 29935 8818 29941 8830
rect 29993 8818 29999 8870
rect 31121 8861 31179 8867
rect 31121 8827 31133 8861
rect 31167 8858 31179 8861
rect 39919 8858 39925 8870
rect 31167 8830 39925 8858
rect 31167 8827 31179 8830
rect 31121 8821 31179 8827
rect 39919 8818 39925 8830
rect 39977 8818 39983 8870
rect 879 7953 939 8009
rect 2127 7953 2187 8009
rect 3375 7953 3435 8009
rect 4623 7953 4683 8009
rect 5871 7953 5931 8009
rect 7119 7953 7179 8009
rect 8367 7953 8427 8009
rect 9615 7953 9675 8009
rect 10863 7953 10923 8009
rect 12111 7953 12171 8009
rect 13359 7953 13419 8009
rect 14607 7953 14667 8009
rect 15855 7953 15915 8009
rect 17103 7953 17163 8009
rect 18351 7953 18411 8009
rect 19599 7953 19659 8009
rect 20847 7953 20907 8009
rect 22095 7953 22155 8009
rect 23343 7953 23403 8009
rect 24591 7953 24651 8009
rect 25839 7953 25899 8009
rect 27087 7953 27147 8009
rect 28335 7953 28395 8009
rect 29583 7953 29643 8009
rect 30831 7953 30891 8009
rect 32079 7953 32139 8009
rect 33327 7953 33387 8009
rect 34575 7953 34635 8009
rect 35823 7953 35883 8009
rect 37071 7953 37131 8009
rect 38319 7953 38379 8009
rect 39567 7953 39627 8009
rect 9967 7919 9973 7928
rect 723 7885 9973 7919
rect 9967 7876 9973 7885
rect 10025 7919 10031 7928
rect 19951 7919 19957 7928
rect 10025 7885 10083 7919
rect 10707 7885 19957 7919
rect 10025 7876 10031 7885
rect 19951 7876 19957 7885
rect 20009 7919 20015 7928
rect 29935 7919 29941 7928
rect 20009 7885 20067 7919
rect 20691 7885 29941 7919
rect 20009 7876 20015 7885
rect 29935 7876 29941 7885
rect 29993 7919 29999 7928
rect 39919 7919 39925 7928
rect 29993 7885 30051 7919
rect 30675 7885 39925 7919
rect 29993 7876 29999 7885
rect 39919 7876 39925 7885
rect 39977 7919 39983 7928
rect 39977 7885 40035 7919
rect 39977 7876 39983 7885
rect 751 5936 779 6002
rect 751 5908 851 5936
rect 728 5496 774 5750
rect 823 4620 851 5908
rect 953 5856 981 6002
rect 1999 5936 2027 6002
rect 1999 5908 2099 5936
rect 896 5828 981 5856
rect 896 4608 924 5828
rect 1976 5496 2022 5750
rect 2071 4620 2099 5908
rect 2201 5856 2229 6002
rect 3247 5936 3275 6002
rect 3247 5908 3347 5936
rect 2144 5828 2229 5856
rect 2144 4608 2172 5828
rect 3224 5496 3270 5750
rect 3319 4620 3347 5908
rect 3449 5856 3477 6002
rect 4495 5936 4523 6002
rect 4495 5908 4595 5936
rect 3392 5828 3477 5856
rect 3392 4608 3420 5828
rect 4472 5496 4518 5750
rect 4567 4620 4595 5908
rect 4697 5856 4725 6002
rect 5743 5936 5771 6002
rect 5743 5908 5843 5936
rect 4640 5828 4725 5856
rect 4640 4608 4668 5828
rect 5720 5496 5766 5750
rect 5815 4620 5843 5908
rect 5945 5856 5973 6002
rect 6991 5936 7019 6002
rect 6991 5908 7091 5936
rect 5888 5828 5973 5856
rect 5888 4608 5916 5828
rect 6968 5496 7014 5750
rect 7063 4620 7091 5908
rect 7193 5856 7221 6002
rect 8239 5936 8267 6002
rect 8239 5908 8339 5936
rect 7136 5828 7221 5856
rect 7136 4608 7164 5828
rect 8216 5496 8262 5750
rect 8311 4620 8339 5908
rect 8441 5856 8469 6002
rect 9487 5936 9515 6002
rect 9487 5908 9587 5936
rect 8384 5828 8469 5856
rect 8384 4608 8412 5828
rect 9464 5496 9510 5750
rect 9559 4620 9587 5908
rect 9689 5856 9717 6002
rect 10735 5936 10763 6002
rect 10735 5908 10835 5936
rect 9632 5828 9717 5856
rect 9632 4608 9660 5828
rect 10712 5496 10758 5750
rect 10807 4620 10835 5908
rect 10937 5856 10965 6002
rect 11983 5936 12011 6002
rect 11983 5908 12083 5936
rect 10880 5828 10965 5856
rect 10880 4608 10908 5828
rect 11960 5496 12006 5750
rect 12055 4620 12083 5908
rect 12185 5856 12213 6002
rect 13231 5936 13259 6002
rect 13231 5908 13331 5936
rect 12128 5828 12213 5856
rect 12128 4608 12156 5828
rect 13208 5496 13254 5750
rect 13303 4620 13331 5908
rect 13433 5856 13461 6002
rect 14479 5936 14507 6002
rect 14479 5908 14579 5936
rect 13376 5828 13461 5856
rect 13376 4608 13404 5828
rect 14456 5496 14502 5750
rect 14551 4620 14579 5908
rect 14681 5856 14709 6002
rect 15727 5936 15755 6002
rect 15727 5908 15827 5936
rect 14624 5828 14709 5856
rect 14624 4608 14652 5828
rect 15704 5496 15750 5750
rect 15799 4620 15827 5908
rect 15929 5856 15957 6002
rect 16975 5936 17003 6002
rect 16975 5908 17075 5936
rect 15872 5828 15957 5856
rect 15872 4608 15900 5828
rect 16952 5496 16998 5750
rect 17047 4620 17075 5908
rect 17177 5856 17205 6002
rect 18223 5936 18251 6002
rect 18223 5908 18323 5936
rect 17120 5828 17205 5856
rect 17120 4608 17148 5828
rect 18200 5496 18246 5750
rect 18295 4620 18323 5908
rect 18425 5856 18453 6002
rect 19471 5936 19499 6002
rect 19471 5908 19571 5936
rect 18368 5828 18453 5856
rect 18368 4608 18396 5828
rect 19448 5496 19494 5750
rect 19543 4620 19571 5908
rect 19673 5856 19701 6002
rect 20719 5936 20747 6002
rect 20719 5908 20819 5936
rect 19616 5828 19701 5856
rect 19616 4608 19644 5828
rect 20696 5496 20742 5750
rect 20791 4620 20819 5908
rect 20921 5856 20949 6002
rect 21967 5936 21995 6002
rect 21967 5908 22067 5936
rect 20864 5828 20949 5856
rect 20864 4608 20892 5828
rect 21944 5496 21990 5750
rect 22039 4620 22067 5908
rect 22169 5856 22197 6002
rect 23215 5936 23243 6002
rect 23215 5908 23315 5936
rect 22112 5828 22197 5856
rect 22112 4608 22140 5828
rect 23192 5496 23238 5750
rect 23287 4620 23315 5908
rect 23417 5856 23445 6002
rect 24463 5936 24491 6002
rect 24463 5908 24563 5936
rect 23360 5828 23445 5856
rect 23360 4608 23388 5828
rect 24440 5496 24486 5750
rect 24535 4620 24563 5908
rect 24665 5856 24693 6002
rect 25711 5936 25739 6002
rect 25711 5908 25811 5936
rect 24608 5828 24693 5856
rect 24608 4608 24636 5828
rect 25688 5496 25734 5750
rect 25783 4620 25811 5908
rect 25913 5856 25941 6002
rect 26959 5936 26987 6002
rect 26959 5908 27059 5936
rect 25856 5828 25941 5856
rect 25856 4608 25884 5828
rect 26936 5496 26982 5750
rect 27031 4620 27059 5908
rect 27161 5856 27189 6002
rect 28207 5936 28235 6002
rect 28207 5908 28307 5936
rect 27104 5828 27189 5856
rect 27104 4608 27132 5828
rect 28184 5496 28230 5750
rect 28279 4620 28307 5908
rect 28409 5856 28437 6002
rect 29455 5936 29483 6002
rect 29455 5908 29555 5936
rect 28352 5828 28437 5856
rect 28352 4608 28380 5828
rect 29432 5496 29478 5750
rect 29527 4620 29555 5908
rect 29657 5856 29685 6002
rect 30703 5936 30731 6002
rect 30703 5908 30803 5936
rect 29600 5828 29685 5856
rect 29600 4608 29628 5828
rect 30680 5496 30726 5750
rect 30775 4620 30803 5908
rect 30905 5856 30933 6002
rect 31951 5936 31979 6002
rect 31951 5908 32051 5936
rect 30848 5828 30933 5856
rect 30848 4608 30876 5828
rect 31928 5496 31974 5750
rect 32023 4620 32051 5908
rect 32153 5856 32181 6002
rect 33199 5936 33227 6002
rect 33199 5908 33299 5936
rect 32096 5828 32181 5856
rect 32096 4608 32124 5828
rect 33176 5496 33222 5750
rect 33271 4620 33299 5908
rect 33401 5856 33429 6002
rect 34447 5936 34475 6002
rect 34447 5908 34547 5936
rect 33344 5828 33429 5856
rect 33344 4608 33372 5828
rect 34424 5496 34470 5750
rect 34519 4620 34547 5908
rect 34649 5856 34677 6002
rect 35695 5936 35723 6002
rect 35695 5908 35795 5936
rect 34592 5828 34677 5856
rect 34592 4608 34620 5828
rect 35672 5496 35718 5750
rect 35767 4620 35795 5908
rect 35897 5856 35925 6002
rect 36943 5936 36971 6002
rect 36943 5908 37043 5936
rect 35840 5828 35925 5856
rect 35840 4608 35868 5828
rect 36920 5496 36966 5750
rect 37015 4620 37043 5908
rect 37145 5856 37173 6002
rect 38191 5936 38219 6002
rect 38191 5908 38291 5936
rect 37088 5828 37173 5856
rect 37088 4608 37116 5828
rect 38168 5496 38214 5750
rect 38263 4620 38291 5908
rect 38393 5856 38421 6002
rect 39439 5936 39467 6002
rect 39439 5908 39539 5936
rect 38336 5828 38421 5856
rect 38336 4608 38364 5828
rect 39416 5496 39462 5750
rect 39511 4620 39539 5908
rect 39641 5856 39669 6002
rect 39584 5828 39669 5856
rect 39584 4608 39612 5828
rect 823 3428 851 3494
rect 704 3400 851 3428
rect 704 2994 732 3400
rect 896 3348 924 3494
rect 2071 3428 2099 3494
rect 1952 3400 2099 3428
rect 896 3320 1196 3348
rect 1168 3118 1196 3320
rect 1952 2994 1980 3400
rect 2144 3348 2172 3494
rect 3319 3428 3347 3494
rect 3200 3400 3347 3428
rect 2144 3320 2444 3348
rect 2416 3118 2444 3320
rect 3200 2994 3228 3400
rect 3392 3348 3420 3494
rect 4567 3428 4595 3494
rect 4448 3400 4595 3428
rect 3392 3320 3692 3348
rect 3664 3118 3692 3320
rect 4448 2994 4476 3400
rect 4640 3348 4668 3494
rect 5815 3428 5843 3494
rect 5696 3400 5843 3428
rect 4640 3320 4940 3348
rect 4912 3118 4940 3320
rect 5696 2994 5724 3400
rect 5888 3348 5916 3494
rect 7063 3428 7091 3494
rect 6944 3400 7091 3428
rect 5888 3320 6188 3348
rect 6160 3118 6188 3320
rect 6944 2994 6972 3400
rect 7136 3348 7164 3494
rect 8311 3428 8339 3494
rect 8192 3400 8339 3428
rect 7136 3320 7436 3348
rect 7408 3118 7436 3320
rect 8192 2994 8220 3400
rect 8384 3348 8412 3494
rect 9559 3428 9587 3494
rect 9440 3400 9587 3428
rect 8384 3320 8684 3348
rect 8656 3118 8684 3320
rect 9440 2994 9468 3400
rect 9632 3348 9660 3494
rect 10807 3428 10835 3494
rect 10688 3400 10835 3428
rect 9632 3320 9932 3348
rect 9904 3118 9932 3320
rect 10688 2994 10716 3400
rect 10880 3348 10908 3494
rect 12055 3428 12083 3494
rect 11936 3400 12083 3428
rect 10880 3320 11180 3348
rect 11152 3118 11180 3320
rect 11936 2994 11964 3400
rect 12128 3348 12156 3494
rect 13303 3428 13331 3494
rect 13184 3400 13331 3428
rect 12128 3320 12428 3348
rect 12400 3118 12428 3320
rect 13184 2994 13212 3400
rect 13376 3348 13404 3494
rect 14551 3428 14579 3494
rect 14432 3400 14579 3428
rect 13376 3320 13676 3348
rect 13648 3118 13676 3320
rect 14432 2994 14460 3400
rect 14624 3348 14652 3494
rect 15799 3428 15827 3494
rect 15680 3400 15827 3428
rect 14624 3320 14924 3348
rect 14896 3118 14924 3320
rect 15680 2994 15708 3400
rect 15872 3348 15900 3494
rect 17047 3428 17075 3494
rect 16928 3400 17075 3428
rect 15872 3320 16172 3348
rect 16144 3118 16172 3320
rect 16928 2994 16956 3400
rect 17120 3348 17148 3494
rect 18295 3428 18323 3494
rect 18176 3400 18323 3428
rect 17120 3320 17420 3348
rect 17392 3118 17420 3320
rect 18176 2994 18204 3400
rect 18368 3348 18396 3494
rect 19543 3428 19571 3494
rect 19424 3400 19571 3428
rect 18368 3320 18668 3348
rect 18640 3118 18668 3320
rect 19424 2994 19452 3400
rect 19616 3348 19644 3494
rect 20791 3428 20819 3494
rect 20672 3400 20819 3428
rect 19616 3320 19916 3348
rect 19888 3118 19916 3320
rect 20672 2994 20700 3400
rect 20864 3348 20892 3494
rect 22039 3428 22067 3494
rect 21920 3400 22067 3428
rect 20864 3320 21164 3348
rect 21136 3118 21164 3320
rect 21920 2994 21948 3400
rect 22112 3348 22140 3494
rect 23287 3428 23315 3494
rect 23168 3400 23315 3428
rect 22112 3320 22412 3348
rect 22384 3118 22412 3320
rect 23168 2994 23196 3400
rect 23360 3348 23388 3494
rect 24535 3428 24563 3494
rect 24416 3400 24563 3428
rect 23360 3320 23660 3348
rect 23632 3118 23660 3320
rect 24416 2994 24444 3400
rect 24608 3348 24636 3494
rect 25783 3428 25811 3494
rect 25664 3400 25811 3428
rect 24608 3320 24908 3348
rect 24880 3118 24908 3320
rect 25664 2994 25692 3400
rect 25856 3348 25884 3494
rect 27031 3428 27059 3494
rect 26912 3400 27059 3428
rect 25856 3320 26156 3348
rect 26128 3118 26156 3320
rect 26912 2994 26940 3400
rect 27104 3348 27132 3494
rect 28279 3428 28307 3494
rect 28160 3400 28307 3428
rect 27104 3320 27404 3348
rect 27376 3118 27404 3320
rect 28160 2994 28188 3400
rect 28352 3348 28380 3494
rect 29527 3428 29555 3494
rect 29408 3400 29555 3428
rect 28352 3320 28652 3348
rect 28624 3118 28652 3320
rect 29408 2994 29436 3400
rect 29600 3348 29628 3494
rect 30775 3428 30803 3494
rect 30656 3400 30803 3428
rect 29600 3320 29900 3348
rect 29872 3118 29900 3320
rect 30656 2994 30684 3400
rect 30848 3348 30876 3494
rect 32023 3428 32051 3494
rect 31904 3400 32051 3428
rect 30848 3320 31148 3348
rect 31120 3118 31148 3320
rect 31904 2994 31932 3400
rect 32096 3348 32124 3494
rect 33271 3428 33299 3494
rect 33152 3400 33299 3428
rect 32096 3320 32396 3348
rect 32368 3118 32396 3320
rect 33152 2994 33180 3400
rect 33344 3348 33372 3494
rect 34519 3428 34547 3494
rect 34400 3400 34547 3428
rect 33344 3320 33644 3348
rect 33616 3118 33644 3320
rect 34400 2994 34428 3400
rect 34592 3348 34620 3494
rect 35767 3428 35795 3494
rect 35648 3400 35795 3428
rect 34592 3320 34892 3348
rect 34864 3118 34892 3320
rect 35648 2994 35676 3400
rect 35840 3348 35868 3494
rect 37015 3428 37043 3494
rect 36896 3400 37043 3428
rect 35840 3320 36140 3348
rect 36112 3118 36140 3320
rect 36896 2994 36924 3400
rect 37088 3348 37116 3494
rect 38263 3428 38291 3494
rect 38144 3400 38291 3428
rect 37088 3320 37388 3348
rect 37360 3118 37388 3320
rect 38144 2994 38172 3400
rect 38336 3348 38364 3494
rect 39511 3428 39539 3494
rect 39392 3400 39539 3428
rect 38336 3320 38636 3348
rect 38608 3118 38636 3320
rect 39392 2994 39420 3400
rect 39584 3348 39612 3494
rect 39584 3320 39884 3348
rect 39856 3118 39884 3320
rect 704 1192 732 1258
rect 690 1164 732 1192
rect 66 252 94 1006
rect 530 252 558 1006
rect 690 252 718 1164
rect 1168 1112 1196 1258
rect 1154 1084 1196 1112
rect 1300 1112 1328 1258
rect 1764 1192 1792 1258
rect 1952 1192 1980 1258
rect 1764 1164 1806 1192
rect 1300 1084 1342 1112
rect 1154 252 1182 1084
rect 1314 252 1342 1084
rect 1778 252 1806 1164
rect 1938 1164 1980 1192
rect 1938 252 1966 1164
rect 2416 1112 2444 1258
rect 2402 1084 2444 1112
rect 2548 1112 2576 1258
rect 3012 1192 3040 1258
rect 3200 1192 3228 1258
rect 3012 1164 3054 1192
rect 2548 1084 2590 1112
rect 2402 252 2430 1084
rect 2562 252 2590 1084
rect 3026 252 3054 1164
rect 3186 1164 3228 1192
rect 3186 252 3214 1164
rect 3664 1112 3692 1258
rect 3650 1084 3692 1112
rect 3796 1112 3824 1258
rect 4260 1192 4288 1258
rect 4448 1192 4476 1258
rect 4260 1164 4302 1192
rect 3796 1084 3838 1112
rect 3650 252 3678 1084
rect 3810 252 3838 1084
rect 4274 252 4302 1164
rect 4434 1164 4476 1192
rect 4434 252 4462 1164
rect 4912 1112 4940 1258
rect 4898 1084 4940 1112
rect 5044 1112 5072 1258
rect 5508 1192 5536 1258
rect 5696 1192 5724 1258
rect 5508 1164 5550 1192
rect 5044 1084 5086 1112
rect 4898 252 4926 1084
rect 5058 252 5086 1084
rect 5522 252 5550 1164
rect 5682 1164 5724 1192
rect 5682 252 5710 1164
rect 6160 1112 6188 1258
rect 6146 1084 6188 1112
rect 6292 1112 6320 1258
rect 6756 1192 6784 1258
rect 6944 1192 6972 1258
rect 6756 1164 6798 1192
rect 6292 1084 6334 1112
rect 6146 252 6174 1084
rect 6306 252 6334 1084
rect 6770 252 6798 1164
rect 6930 1164 6972 1192
rect 6930 252 6958 1164
rect 7408 1112 7436 1258
rect 7394 1084 7436 1112
rect 7540 1112 7568 1258
rect 8004 1192 8032 1258
rect 8192 1192 8220 1258
rect 8004 1164 8046 1192
rect 7540 1084 7582 1112
rect 7394 252 7422 1084
rect 7554 252 7582 1084
rect 8018 252 8046 1164
rect 8178 1164 8220 1192
rect 8178 252 8206 1164
rect 8656 1112 8684 1258
rect 8642 1084 8684 1112
rect 8788 1112 8816 1258
rect 9252 1192 9280 1258
rect 9440 1192 9468 1258
rect 9252 1164 9294 1192
rect 8788 1084 8830 1112
rect 8642 252 8670 1084
rect 8802 252 8830 1084
rect 9266 252 9294 1164
rect 9426 1164 9468 1192
rect 9426 252 9454 1164
rect 9904 1112 9932 1258
rect 9890 1084 9932 1112
rect 10036 1112 10064 1258
rect 10500 1192 10528 1258
rect 10688 1192 10716 1258
rect 10500 1164 10542 1192
rect 10036 1084 10078 1112
rect 9890 252 9918 1084
rect 10050 252 10078 1084
rect 10514 252 10542 1164
rect 10674 1164 10716 1192
rect 10674 252 10702 1164
rect 11152 1112 11180 1258
rect 11138 1084 11180 1112
rect 11284 1112 11312 1258
rect 11748 1192 11776 1258
rect 11936 1192 11964 1258
rect 11748 1164 11790 1192
rect 11284 1084 11326 1112
rect 11138 252 11166 1084
rect 11298 252 11326 1084
rect 11762 252 11790 1164
rect 11922 1164 11964 1192
rect 11922 252 11950 1164
rect 12400 1112 12428 1258
rect 12386 1084 12428 1112
rect 12532 1112 12560 1258
rect 12996 1192 13024 1258
rect 13184 1192 13212 1258
rect 12996 1164 13038 1192
rect 12532 1084 12574 1112
rect 12386 252 12414 1084
rect 12546 252 12574 1084
rect 13010 252 13038 1164
rect 13170 1164 13212 1192
rect 13170 252 13198 1164
rect 13648 1112 13676 1258
rect 13634 1084 13676 1112
rect 13780 1112 13808 1258
rect 14244 1192 14272 1258
rect 14432 1192 14460 1258
rect 14244 1164 14286 1192
rect 13780 1084 13822 1112
rect 13634 252 13662 1084
rect 13794 252 13822 1084
rect 14258 252 14286 1164
rect 14418 1164 14460 1192
rect 14418 252 14446 1164
rect 14896 1112 14924 1258
rect 14882 1084 14924 1112
rect 15028 1112 15056 1258
rect 15492 1192 15520 1258
rect 15680 1192 15708 1258
rect 15492 1164 15534 1192
rect 15028 1084 15070 1112
rect 14882 252 14910 1084
rect 15042 252 15070 1084
rect 15506 252 15534 1164
rect 15666 1164 15708 1192
rect 15666 252 15694 1164
rect 16144 1112 16172 1258
rect 16130 1084 16172 1112
rect 16276 1112 16304 1258
rect 16740 1192 16768 1258
rect 16928 1192 16956 1258
rect 16740 1164 16782 1192
rect 16276 1084 16318 1112
rect 16130 252 16158 1084
rect 16290 252 16318 1084
rect 16754 252 16782 1164
rect 16914 1164 16956 1192
rect 16914 252 16942 1164
rect 17392 1112 17420 1258
rect 17378 1084 17420 1112
rect 17524 1112 17552 1258
rect 17988 1192 18016 1258
rect 18176 1192 18204 1258
rect 17988 1164 18030 1192
rect 17524 1084 17566 1112
rect 17378 252 17406 1084
rect 17538 252 17566 1084
rect 18002 252 18030 1164
rect 18162 1164 18204 1192
rect 18162 252 18190 1164
rect 18640 1112 18668 1258
rect 18626 1084 18668 1112
rect 18772 1112 18800 1258
rect 19236 1192 19264 1258
rect 19424 1192 19452 1258
rect 19236 1164 19278 1192
rect 18772 1084 18814 1112
rect 18626 252 18654 1084
rect 18786 252 18814 1084
rect 19250 252 19278 1164
rect 19410 1164 19452 1192
rect 19410 252 19438 1164
rect 19888 1112 19916 1258
rect 19874 1084 19916 1112
rect 20020 1112 20048 1258
rect 20484 1192 20512 1258
rect 20672 1192 20700 1258
rect 20484 1164 20526 1192
rect 20020 1084 20062 1112
rect 19874 252 19902 1084
rect 20034 252 20062 1084
rect 20498 252 20526 1164
rect 20658 1164 20700 1192
rect 20658 252 20686 1164
rect 21136 1112 21164 1258
rect 21122 1084 21164 1112
rect 21268 1112 21296 1258
rect 21732 1192 21760 1258
rect 21920 1192 21948 1258
rect 21732 1164 21774 1192
rect 21268 1084 21310 1112
rect 21122 252 21150 1084
rect 21282 252 21310 1084
rect 21746 252 21774 1164
rect 21906 1164 21948 1192
rect 21906 252 21934 1164
rect 22384 1112 22412 1258
rect 22370 1084 22412 1112
rect 22516 1112 22544 1258
rect 22980 1192 23008 1258
rect 23168 1192 23196 1258
rect 22980 1164 23022 1192
rect 22516 1084 22558 1112
rect 22370 252 22398 1084
rect 22530 252 22558 1084
rect 22994 252 23022 1164
rect 23154 1164 23196 1192
rect 23154 252 23182 1164
rect 23632 1112 23660 1258
rect 23618 1084 23660 1112
rect 23764 1112 23792 1258
rect 24228 1192 24256 1258
rect 24416 1192 24444 1258
rect 24228 1164 24270 1192
rect 23764 1084 23806 1112
rect 23618 252 23646 1084
rect 23778 252 23806 1084
rect 24242 252 24270 1164
rect 24402 1164 24444 1192
rect 24402 252 24430 1164
rect 24880 1112 24908 1258
rect 24866 1084 24908 1112
rect 25012 1112 25040 1258
rect 25476 1192 25504 1258
rect 25664 1192 25692 1258
rect 25476 1164 25518 1192
rect 25012 1084 25054 1112
rect 24866 252 24894 1084
rect 25026 252 25054 1084
rect 25490 252 25518 1164
rect 25650 1164 25692 1192
rect 25650 252 25678 1164
rect 26128 1112 26156 1258
rect 26114 1084 26156 1112
rect 26260 1112 26288 1258
rect 26724 1192 26752 1258
rect 26912 1192 26940 1258
rect 26724 1164 26766 1192
rect 26260 1084 26302 1112
rect 26114 252 26142 1084
rect 26274 252 26302 1084
rect 26738 252 26766 1164
rect 26898 1164 26940 1192
rect 26898 252 26926 1164
rect 27376 1112 27404 1258
rect 27362 1084 27404 1112
rect 27508 1112 27536 1258
rect 27972 1192 28000 1258
rect 28160 1192 28188 1258
rect 27972 1164 28014 1192
rect 27508 1084 27550 1112
rect 27362 252 27390 1084
rect 27522 252 27550 1084
rect 27986 252 28014 1164
rect 28146 1164 28188 1192
rect 28146 252 28174 1164
rect 28624 1112 28652 1258
rect 28610 1084 28652 1112
rect 28756 1112 28784 1258
rect 29220 1192 29248 1258
rect 29408 1192 29436 1258
rect 29220 1164 29262 1192
rect 28756 1084 28798 1112
rect 28610 252 28638 1084
rect 28770 252 28798 1084
rect 29234 252 29262 1164
rect 29394 1164 29436 1192
rect 29394 252 29422 1164
rect 29872 1112 29900 1258
rect 29858 1084 29900 1112
rect 30004 1112 30032 1258
rect 30468 1192 30496 1258
rect 30656 1192 30684 1258
rect 30468 1164 30510 1192
rect 30004 1084 30046 1112
rect 29858 252 29886 1084
rect 30018 252 30046 1084
rect 30482 252 30510 1164
rect 30642 1164 30684 1192
rect 30642 252 30670 1164
rect 31120 1112 31148 1258
rect 31106 1084 31148 1112
rect 31252 1112 31280 1258
rect 31716 1192 31744 1258
rect 31904 1192 31932 1258
rect 31716 1164 31758 1192
rect 31252 1084 31294 1112
rect 31106 252 31134 1084
rect 31266 252 31294 1084
rect 31730 252 31758 1164
rect 31890 1164 31932 1192
rect 31890 252 31918 1164
rect 32368 1112 32396 1258
rect 32354 1084 32396 1112
rect 32500 1112 32528 1258
rect 32964 1192 32992 1258
rect 33152 1192 33180 1258
rect 32964 1164 33006 1192
rect 32500 1084 32542 1112
rect 32354 252 32382 1084
rect 32514 252 32542 1084
rect 32978 252 33006 1164
rect 33138 1164 33180 1192
rect 33138 252 33166 1164
rect 33616 1112 33644 1258
rect 33602 1084 33644 1112
rect 33748 1112 33776 1258
rect 34212 1192 34240 1258
rect 34400 1192 34428 1258
rect 34212 1164 34254 1192
rect 33748 1084 33790 1112
rect 33602 252 33630 1084
rect 33762 252 33790 1084
rect 34226 252 34254 1164
rect 34386 1164 34428 1192
rect 34386 252 34414 1164
rect 34864 1112 34892 1258
rect 34850 1084 34892 1112
rect 34996 1112 35024 1258
rect 35460 1192 35488 1258
rect 35648 1192 35676 1258
rect 35460 1164 35502 1192
rect 34996 1084 35038 1112
rect 34850 252 34878 1084
rect 35010 252 35038 1084
rect 35474 252 35502 1164
rect 35634 1164 35676 1192
rect 35634 252 35662 1164
rect 36112 1112 36140 1258
rect 36098 1084 36140 1112
rect 36244 1112 36272 1258
rect 36708 1192 36736 1258
rect 36896 1192 36924 1258
rect 36708 1164 36750 1192
rect 36244 1084 36286 1112
rect 36098 252 36126 1084
rect 36258 252 36286 1084
rect 36722 252 36750 1164
rect 36882 1164 36924 1192
rect 36882 252 36910 1164
rect 37360 1112 37388 1258
rect 37346 1084 37388 1112
rect 37492 1112 37520 1258
rect 37956 1192 37984 1258
rect 38144 1192 38172 1258
rect 37956 1164 37998 1192
rect 37492 1084 37534 1112
rect 37346 252 37374 1084
rect 37506 252 37534 1084
rect 37970 252 37998 1164
rect 38130 1164 38172 1192
rect 38130 252 38158 1164
rect 38608 1112 38636 1258
rect 38594 1084 38636 1112
rect 38740 1112 38768 1258
rect 39204 1192 39232 1258
rect 39392 1192 39420 1258
rect 39204 1164 39246 1192
rect 38740 1084 38782 1112
rect 38594 252 38622 1084
rect 38754 252 38782 1084
rect 39218 252 39246 1164
rect 39378 1164 39420 1192
rect 39378 252 39406 1164
rect 39856 1112 39884 1258
rect 39842 1084 39884 1112
rect 39988 1112 40016 1258
rect 40452 1192 40480 1258
rect 40452 1164 40494 1192
rect 39988 1084 40030 1112
rect 39842 252 39870 1084
rect 40002 252 40030 1084
rect 40466 252 40494 1164
<< via1 >>
rect 9973 8818 10025 8870
rect 19957 8818 20009 8870
rect 29941 8818 29993 8870
rect 39925 8818 39977 8870
rect 9973 7876 10025 7928
rect 19957 7876 20009 7928
rect 29941 7876 29993 7928
rect 39925 7876 39977 7928
<< metal2 >>
rect 610 9101 638 9129
rect 10594 9101 10622 9129
rect 20578 9101 20606 9129
rect 30562 9101 30590 9129
rect 9973 8870 10025 8876
rect 9973 8812 10025 8818
rect 19957 8870 20009 8876
rect 19957 8812 20009 8818
rect 29941 8870 29993 8876
rect 29941 8812 29993 8818
rect 39925 8870 39977 8876
rect 39925 8812 39977 8818
rect 9985 7934 10013 8812
rect 19969 7934 19997 8812
rect 29953 7934 29981 8812
rect 39937 7934 39965 8812
rect 9973 7928 10025 7934
rect 9973 7870 10025 7876
rect 19957 7928 20009 7934
rect 19957 7870 20009 7876
rect 29941 7928 29993 7934
rect 29941 7870 29993 7876
rect 39925 7928 39977 7934
rect 39925 7870 39977 7876
<< metal3 >>
rect 948 9336 1046 9434
rect 10932 9336 11030 9434
rect 20916 9336 21014 9434
rect 30900 9336 30998 9434
rect 624 8837 40560 8897
rect 948 8216 1046 8314
rect 10932 8216 11030 8314
rect 20916 8216 21014 8314
rect 30900 8216 30998 8314
rect 851 7773 949 7871
rect 2099 7773 2197 7871
rect 3347 7773 3445 7871
rect 4595 7773 4693 7871
rect 5843 7773 5941 7871
rect 7091 7773 7189 7871
rect 8339 7773 8437 7871
rect 9587 7773 9685 7871
rect 10835 7773 10933 7871
rect 12083 7773 12181 7871
rect 13331 7773 13429 7871
rect 14579 7773 14677 7871
rect 15827 7773 15925 7871
rect 17075 7773 17173 7871
rect 18323 7773 18421 7871
rect 19571 7773 19669 7871
rect 20819 7773 20917 7871
rect 22067 7773 22165 7871
rect 23315 7773 23413 7871
rect 24563 7773 24661 7871
rect 25811 7773 25909 7871
rect 27059 7773 27157 7871
rect 28307 7773 28405 7871
rect 29555 7773 29653 7871
rect 30803 7773 30901 7871
rect 32051 7773 32149 7871
rect 33299 7773 33397 7871
rect 34547 7773 34645 7871
rect 35795 7773 35893 7871
rect 37043 7773 37141 7871
rect 38291 7773 38389 7871
rect 39539 7773 39637 7871
rect 837 7357 935 7455
rect 2085 7357 2183 7455
rect 3333 7357 3431 7455
rect 4581 7357 4679 7455
rect 5829 7357 5927 7455
rect 7077 7357 7175 7455
rect 8325 7357 8423 7455
rect 9573 7357 9671 7455
rect 10821 7357 10919 7455
rect 12069 7357 12167 7455
rect 13317 7357 13415 7455
rect 14565 7357 14663 7455
rect 15813 7357 15911 7455
rect 17061 7357 17159 7455
rect 18309 7357 18407 7455
rect 19557 7357 19655 7455
rect 20805 7357 20903 7455
rect 22053 7357 22151 7455
rect 23301 7357 23399 7455
rect 24549 7357 24647 7455
rect 25797 7357 25895 7455
rect 27045 7357 27143 7455
rect 28293 7357 28391 7455
rect 29541 7357 29639 7455
rect 30789 7357 30887 7455
rect 32037 7357 32135 7455
rect 33285 7357 33383 7455
rect 34533 7357 34631 7455
rect 35781 7357 35879 7455
rect 37029 7357 37127 7455
rect 38277 7357 38375 7455
rect 39525 7357 39623 7455
rect 952 7155 1050 7253
rect 2200 7155 2298 7253
rect 3448 7155 3546 7253
rect 4696 7155 4794 7253
rect 5944 7155 6042 7253
rect 7192 7155 7290 7253
rect 8440 7155 8538 7253
rect 9688 7155 9786 7253
rect 10936 7155 11034 7253
rect 12184 7155 12282 7253
rect 13432 7155 13530 7253
rect 14680 7155 14778 7253
rect 15928 7155 16026 7253
rect 17176 7155 17274 7253
rect 18424 7155 18522 7253
rect 19672 7155 19770 7253
rect 20920 7155 21018 7253
rect 22168 7155 22266 7253
rect 23416 7155 23514 7253
rect 24664 7155 24762 7253
rect 25912 7155 26010 7253
rect 27160 7155 27258 7253
rect 28408 7155 28506 7253
rect 29656 7155 29754 7253
rect 30904 7155 31002 7253
rect 32152 7155 32250 7253
rect 33400 7155 33498 7253
rect 34648 7155 34746 7253
rect 35896 7155 35994 7253
rect 37144 7155 37242 7253
rect 38392 7155 38490 7253
rect 39640 7155 39738 7253
rect 831 6823 929 6921
rect 2079 6823 2177 6921
rect 3327 6823 3425 6921
rect 4575 6823 4673 6921
rect 5823 6823 5921 6921
rect 7071 6823 7169 6921
rect 8319 6823 8417 6921
rect 9567 6823 9665 6921
rect 10815 6823 10913 6921
rect 12063 6823 12161 6921
rect 13311 6823 13409 6921
rect 14559 6823 14657 6921
rect 15807 6823 15905 6921
rect 17055 6823 17153 6921
rect 18303 6823 18401 6921
rect 19551 6823 19649 6921
rect 20799 6823 20897 6921
rect 22047 6823 22145 6921
rect 23295 6823 23393 6921
rect 24543 6823 24641 6921
rect 25791 6823 25889 6921
rect 27039 6823 27137 6921
rect 28287 6823 28385 6921
rect 29535 6823 29633 6921
rect 30783 6823 30881 6921
rect 32031 6823 32129 6921
rect 33279 6823 33377 6921
rect 34527 6823 34625 6921
rect 35775 6823 35873 6921
rect 37023 6823 37121 6921
rect 38271 6823 38369 6921
rect 39519 6823 39617 6921
rect 842 6386 940 6484
rect 2090 6386 2188 6484
rect 3338 6386 3436 6484
rect 4586 6386 4684 6484
rect 5834 6386 5932 6484
rect 7082 6386 7180 6484
rect 8330 6386 8428 6484
rect 9578 6386 9676 6484
rect 10826 6386 10924 6484
rect 12074 6386 12172 6484
rect 13322 6386 13420 6484
rect 14570 6386 14668 6484
rect 15818 6386 15916 6484
rect 17066 6386 17164 6484
rect 18314 6386 18412 6484
rect 19562 6386 19660 6484
rect 20810 6386 20908 6484
rect 22058 6386 22156 6484
rect 23306 6386 23404 6484
rect 24554 6386 24652 6484
rect 25802 6386 25900 6484
rect 27050 6386 27148 6484
rect 28298 6386 28396 6484
rect 29546 6386 29644 6484
rect 30794 6386 30892 6484
rect 32042 6386 32140 6484
rect 33290 6386 33388 6484
rect 34538 6386 34636 6484
rect 35786 6386 35884 6484
rect 37034 6386 37132 6484
rect 38282 6386 38380 6484
rect 39530 6386 39628 6484
rect 956 5593 1054 5691
rect 2204 5593 2302 5691
rect 3452 5593 3550 5691
rect 4700 5593 4798 5691
rect 5948 5593 6046 5691
rect 7196 5593 7294 5691
rect 8444 5593 8542 5691
rect 9692 5593 9790 5691
rect 10940 5593 11038 5691
rect 12188 5593 12286 5691
rect 13436 5593 13534 5691
rect 14684 5593 14782 5691
rect 15932 5593 16030 5691
rect 17180 5593 17278 5691
rect 18428 5593 18526 5691
rect 19676 5593 19774 5691
rect 20924 5593 21022 5691
rect 22172 5593 22270 5691
rect 23420 5593 23518 5691
rect 24668 5593 24766 5691
rect 25916 5593 26014 5691
rect 27164 5593 27262 5691
rect 28412 5593 28510 5691
rect 29660 5593 29758 5691
rect 30908 5593 31006 5691
rect 32156 5593 32254 5691
rect 33404 5593 33502 5691
rect 34652 5593 34750 5691
rect 35900 5593 35998 5691
rect 37148 5593 37246 5691
rect 38396 5593 38494 5691
rect 39644 5593 39742 5691
rect 956 5271 1054 5369
rect 2204 5271 2302 5369
rect 3452 5271 3550 5369
rect 4700 5271 4798 5369
rect 5948 5271 6046 5369
rect 7196 5271 7294 5369
rect 8444 5271 8542 5369
rect 9692 5271 9790 5369
rect 10940 5271 11038 5369
rect 12188 5271 12286 5369
rect 13436 5271 13534 5369
rect 14684 5271 14782 5369
rect 15932 5271 16030 5369
rect 17180 5271 17278 5369
rect 18428 5271 18526 5369
rect 19676 5271 19774 5369
rect 20924 5271 21022 5369
rect 22172 5271 22270 5369
rect 23420 5271 23518 5369
rect 24668 5271 24766 5369
rect 25916 5271 26014 5369
rect 27164 5271 27262 5369
rect 28412 5271 28510 5369
rect 29660 5271 29758 5369
rect 30908 5271 31006 5369
rect 32156 5271 32254 5369
rect 33404 5271 33502 5369
rect 34652 5271 34750 5369
rect 35900 5271 35998 5369
rect 37148 5271 37246 5369
rect 38396 5271 38494 5369
rect 39644 5271 39742 5369
rect 944 4433 1042 4531
rect 2192 4433 2290 4531
rect 3440 4433 3538 4531
rect 4688 4433 4786 4531
rect 5936 4433 6034 4531
rect 7184 4433 7282 4531
rect 8432 4433 8530 4531
rect 9680 4433 9778 4531
rect 10928 4433 11026 4531
rect 12176 4433 12274 4531
rect 13424 4433 13522 4531
rect 14672 4433 14770 4531
rect 15920 4433 16018 4531
rect 17168 4433 17266 4531
rect 18416 4433 18514 4531
rect 19664 4433 19762 4531
rect 20912 4433 21010 4531
rect 22160 4433 22258 4531
rect 23408 4433 23506 4531
rect 24656 4433 24754 4531
rect 25904 4433 26002 4531
rect 27152 4433 27250 4531
rect 28400 4433 28498 4531
rect 29648 4433 29746 4531
rect 30896 4433 30994 4531
rect 32144 4433 32242 4531
rect 33392 4433 33490 4531
rect 34640 4433 34738 4531
rect 35888 4433 35986 4531
rect 37136 4433 37234 4531
rect 38384 4433 38482 4531
rect 39632 4433 39730 4531
rect 1026 3659 1124 3757
rect 2274 3659 2372 3757
rect 3522 3659 3620 3757
rect 4770 3659 4868 3757
rect 6018 3659 6116 3757
rect 7266 3659 7364 3757
rect 8514 3659 8612 3757
rect 9762 3659 9860 3757
rect 11010 3659 11108 3757
rect 12258 3659 12356 3757
rect 13506 3659 13604 3757
rect 14754 3659 14852 3757
rect 16002 3659 16100 3757
rect 17250 3659 17348 3757
rect 18498 3659 18596 3757
rect 19746 3659 19844 3757
rect 20994 3659 21092 3757
rect 22242 3659 22340 3757
rect 23490 3659 23588 3757
rect 24738 3659 24836 3757
rect 25986 3659 26084 3757
rect 27234 3659 27332 3757
rect 28482 3659 28580 3757
rect 29730 3659 29828 3757
rect 30978 3659 31076 3757
rect 32226 3659 32324 3757
rect 33474 3659 33572 3757
rect 34722 3659 34820 3757
rect 35970 3659 36068 3757
rect 37218 3659 37316 3757
rect 38466 3659 38564 3757
rect 39714 3659 39812 3757
rect 624 3526 40560 3586
rect 624 2810 40560 2870
rect 624 2686 40560 2746
rect 1199 1886 1297 1984
rect 2447 1886 2545 1984
rect 3695 1886 3793 1984
rect 4943 1886 5041 1984
rect 6191 1886 6289 1984
rect 7439 1886 7537 1984
rect 8687 1886 8785 1984
rect 9935 1886 10033 1984
rect 11183 1886 11281 1984
rect 12431 1886 12529 1984
rect 13679 1886 13777 1984
rect 14927 1886 15025 1984
rect 16175 1886 16273 1984
rect 17423 1886 17521 1984
rect 18671 1886 18769 1984
rect 19919 1886 20017 1984
rect 21167 1886 21265 1984
rect 22415 1886 22513 1984
rect 23663 1886 23761 1984
rect 24911 1886 25009 1984
rect 26159 1886 26257 1984
rect 27407 1886 27505 1984
rect 28655 1886 28753 1984
rect 29903 1886 30001 1984
rect 31151 1886 31249 1984
rect 32399 1886 32497 1984
rect 33647 1886 33745 1984
rect 34895 1886 34993 1984
rect 36143 1886 36241 1984
rect 37391 1886 37489 1984
rect 38639 1886 38737 1984
rect 39887 1886 39985 1984
rect 0 951 40560 1011
rect 382 313 480 411
rect 768 313 866 411
rect 1630 313 1728 411
rect 2016 313 2114 411
rect 2878 313 2976 411
rect 3264 313 3362 411
rect 4126 313 4224 411
rect 4512 313 4610 411
rect 5374 313 5472 411
rect 5760 313 5858 411
rect 6622 313 6720 411
rect 7008 313 7106 411
rect 7870 313 7968 411
rect 8256 313 8354 411
rect 9118 313 9216 411
rect 9504 313 9602 411
rect 10366 313 10464 411
rect 10752 313 10850 411
rect 11614 313 11712 411
rect 12000 313 12098 411
rect 12862 313 12960 411
rect 13248 313 13346 411
rect 14110 313 14208 411
rect 14496 313 14594 411
rect 15358 313 15456 411
rect 15744 313 15842 411
rect 16606 313 16704 411
rect 16992 313 17090 411
rect 17854 313 17952 411
rect 18240 313 18338 411
rect 19102 313 19200 411
rect 19488 313 19586 411
rect 20350 313 20448 411
rect 20736 313 20834 411
rect 21598 313 21696 411
rect 21984 313 22082 411
rect 22846 313 22944 411
rect 23232 313 23330 411
rect 24094 313 24192 411
rect 24480 313 24578 411
rect 25342 313 25440 411
rect 25728 313 25826 411
rect 26590 313 26688 411
rect 26976 313 27074 411
rect 27838 313 27936 411
rect 28224 313 28322 411
rect 29086 313 29184 411
rect 29472 313 29570 411
rect 30334 313 30432 411
rect 30720 313 30818 411
rect 31582 313 31680 411
rect 31968 313 32066 411
rect 32830 313 32928 411
rect 33216 313 33314 411
rect 34078 313 34176 411
rect 34464 313 34562 411
rect 35326 313 35424 411
rect 35712 313 35810 411
rect 36574 313 36672 411
rect 36960 313 37058 411
rect 37822 313 37920 411
rect 38208 313 38306 411
rect 39070 313 39168 411
rect 39456 313 39554 411
rect 40318 313 40416 411
use contact_7  contact_7_0
timestamp 1676037725
transform 1 0 31121 0 1 8811
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1676037725
transform 1 0 21137 0 1 8811
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1676037725
transform 1 0 11153 0 1 8811
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1676037725
transform 1 0 1169 0 1 8811
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1676037725
transform 1 0 39919 0 1 8812
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1676037725
transform 1 0 39919 0 1 7870
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1676037725
transform 1 0 29935 0 1 8812
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1676037725
transform 1 0 29935 0 1 7870
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1676037725
transform 1 0 19951 0 1 8812
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1676037725
transform 1 0 19951 0 1 7870
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1676037725
transform 1 0 9967 0 1 8812
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1676037725
transform 1 0 9967 0 1 7870
box 0 0 1 1
use precharge_array  precharge_array_0
timestamp 1676037725
transform 1 0 0 0 -1 1006
box 0 -12 40560 768
use sense_amp_array  sense_amp_array_0
timestamp 1676037725
transform 1 0 624 0 -1 5750
box -160 0 39936 2256
use single_level_column_mux_array  single_level_column_mux_array_0
timestamp 1676037725
transform 1 0 624 0 -1 3242
box 0 87 39936 1984
use write_driver_array  write_driver_array_0
timestamp 1676037725
transform 1 0 624 0 -1 8013
box -152 4 39411 2011
use write_mask_and_array  write_mask_and_array_0
timestamp 1676037725
transform 1 0 624 0 -1 9385
box -36 -49 39936 1177
<< labels >>
rlabel locali s 11182 8844 11182 8844 4 wdriver_sel_1
port 1 nsew
rlabel locali s 21166 8844 21166 8844 4 wdriver_sel_2
port 2 nsew
rlabel locali s 1198 8844 1198 8844 4 wdriver_sel_0
port 3 nsew
rlabel locali s 31150 8844 31150 8844 4 wdriver_sel_3
port 4 nsew
rlabel metal1 s 29613 7981 29613 7981 4 din_23
port 58 nsew
rlabel metal1 s 26959 5623 26959 5623 4 dout_21
port 24 nsew
rlabel metal1 s 31951 5623 31951 5623 4 dout_25
port 28 nsew
rlabel metal1 s 27117 7981 27117 7981 4 din_21
port 56 nsew
rlabel metal1 s 38191 5623 38191 5623 4 dout_30
port 33 nsew
rlabel metal1 s 34605 7981 34605 7981 4 din_27
port 62 nsew
rlabel metal1 s 30703 5623 30703 5623 4 dout_24
port 27 nsew
rlabel metal1 s 24621 7981 24621 7981 4 din_19
port 54 nsew
rlabel metal1 s 35695 5623 35695 5623 4 dout_28
port 31 nsew
rlabel metal1 s 33199 5623 33199 5623 4 dout_26
port 29 nsew
rlabel metal1 s 30861 7981 30861 7981 4 din_24
port 59 nsew
rlabel metal1 s 23215 5623 23215 5623 4 dout_18
port 21 nsew
rlabel metal1 s 28207 5623 28207 5623 4 dout_22
port 25 nsew
rlabel metal1 s 20719 5623 20719 5623 4 dout_16
port 19 nsew
rlabel metal1 s 23373 7981 23373 7981 4 din_18
port 53 nsew
rlabel metal1 s 36943 5623 36943 5623 4 dout_29
port 32 nsew
rlabel metal1 s 39597 7981 39597 7981 4 din_31
port 66 nsew
rlabel metal1 s 37101 7981 37101 7981 4 din_29
port 64 nsew
rlabel metal1 s 33357 7981 33357 7981 4 din_26
port 61 nsew
rlabel metal1 s 20877 7981 20877 7981 4 din_16
port 51 nsew
rlabel metal1 s 32109 7981 32109 7981 4 din_25
port 60 nsew
rlabel metal1 s 29455 5623 29455 5623 4 dout_23
port 26 nsew
rlabel metal1 s 25371 7902 25371 7902 4 wdriver_sel_2
port 2 nsew
rlabel metal1 s 35853 7981 35853 7981 4 din_28
port 63 nsew
rlabel metal1 s 22125 7981 22125 7981 4 din_17
port 52 nsew
rlabel metal1 s 25869 7981 25869 7981 4 din_20
port 55 nsew
rlabel metal1 s 24463 5623 24463 5623 4 dout_19
port 22 nsew
rlabel metal1 s 39439 5623 39439 5623 4 dout_31
port 34 nsew
rlabel metal1 s 25711 5623 25711 5623 4 dout_20
port 23 nsew
rlabel metal1 s 35355 7902 35355 7902 4 wdriver_sel_3
port 4 nsew
rlabel metal1 s 28365 7981 28365 7981 4 din_22
port 57 nsew
rlabel metal1 s 38349 7981 38349 7981 4 din_30
port 65 nsew
rlabel metal1 s 21967 5623 21967 5623 4 dout_17
port 20 nsew
rlabel metal1 s 34447 5623 34447 5623 4 dout_27
port 30 nsew
rlabel metal1 s 3405 7981 3405 7981 4 din_2
port 37 nsew
rlabel metal1 s 1999 5623 1999 5623 4 dout_1
port 4 nsew
rlabel metal1 s 19629 7981 19629 7981 4 din_15
port 50 nsew
rlabel metal1 s 12141 7981 12141 7981 4 din_9
port 44 nsew
rlabel metal1 s 9645 7981 9645 7981 4 din_7
port 42 nsew
rlabel metal1 s 8397 7981 8397 7981 4 din_6
port 41 nsew
rlabel metal1 s 909 7981 909 7981 4 din_0
port 35 nsew
rlabel metal1 s 17133 7981 17133 7981 4 din_13
port 48 nsew
rlabel metal1 s 5901 7981 5901 7981 4 din_4
port 39 nsew
rlabel metal1 s 6991 5623 6991 5623 4 dout_5
port 8 nsew
rlabel metal1 s 18381 7981 18381 7981 4 din_14
port 49 nsew
rlabel metal1 s 751 5623 751 5623 4 dout_0
port 3 nsew
rlabel metal1 s 5403 7902 5403 7902 4 wdriver_sel_0
port 3 nsew
rlabel metal1 s 4653 7981 4653 7981 4 din_3
port 38 nsew
rlabel metal1 s 13231 5623 13231 5623 4 dout_10
port 13 nsew
rlabel metal1 s 15885 7981 15885 7981 4 din_12
port 47 nsew
rlabel metal1 s 9487 5623 9487 5623 4 dout_7
port 10 nsew
rlabel metal1 s 10893 7981 10893 7981 4 din_8
port 43 nsew
rlabel metal1 s 11983 5623 11983 5623 4 dout_9
port 12 nsew
rlabel metal1 s 19471 5623 19471 5623 4 dout_15
port 18 nsew
rlabel metal1 s 8239 5623 8239 5623 4 dout_6
port 9 nsew
rlabel metal1 s 10735 5623 10735 5623 4 dout_8
port 11 nsew
rlabel metal1 s 15387 7902 15387 7902 4 wdriver_sel_1
port 1 nsew
rlabel metal1 s 4495 5623 4495 5623 4 dout_3
port 6 nsew
rlabel metal1 s 2157 7981 2157 7981 4 din_1
port 36 nsew
rlabel metal1 s 13389 7981 13389 7981 4 din_10
port 45 nsew
rlabel metal1 s 3247 5623 3247 5623 4 dout_2
port 5 nsew
rlabel metal1 s 5743 5623 5743 5623 4 dout_4
port 7 nsew
rlabel metal1 s 14637 7981 14637 7981 4 din_11
port 46 nsew
rlabel metal1 s 16975 5623 16975 5623 4 dout_13
port 16 nsew
rlabel metal1 s 14479 5623 14479 5623 4 dout_11
port 14 nsew
rlabel metal1 s 18223 5623 18223 5623 4 dout_14
port 17 nsew
rlabel metal1 s 7149 7981 7149 7981 4 din_5
port 40 nsew
rlabel metal1 s 15727 5623 15727 5623 4 dout_12
port 15 nsew
rlabel metal1 s 10688 629 10688 629 4 bl_16
port 35 nsew
rlabel metal1 s 15520 629 15520 629 4 bl_23
port 49 nsew
rlabel metal1 s 7568 629 7568 629 4 br_11
port 26 nsew
rlabel metal1 s 1952 629 1952 629 4 bl_2
port 7 nsew
rlabel metal1 s 8656 629 8656 629 4 br_12
port 28 nsew
rlabel metal1 s 19424 629 19424 629 4 bl_30
port 63 nsew
rlabel metal1 s 15056 629 15056 629 4 br_23
port 50 nsew
rlabel metal1 s 1328 629 1328 629 4 br_1
port 6 nsew
rlabel metal1 s 12400 629 12400 629 4 br_18
port 40 nsew
rlabel metal1 s 1792 629 1792 629 4 bl_1
port 5 nsew
rlabel metal1 s 17392 629 17392 629 4 br_26
port 56 nsew
rlabel metal1 s 11312 629 11312 629 4 br_17
port 38 nsew
rlabel metal1 s 16928 629 16928 629 4 bl_26
port 55 nsew
rlabel metal1 s 13184 629 13184 629 4 bl_20
port 43 nsew
rlabel metal1 s 5536 629 5536 629 4 bl_7
port 17 nsew
rlabel metal1 s 11776 629 11776 629 4 bl_17
port 37 nsew
rlabel metal1 s 3040 629 3040 629 4 bl_3
port 9 nsew
rlabel metal1 s 13808 629 13808 629 4 br_21
port 46 nsew
rlabel metal1 s 11936 629 11936 629 4 bl_18
port 39 nsew
rlabel metal1 s 8192 629 8192 629 4 bl_12
port 27 nsew
rlabel metal1 s 8816 629 8816 629 4 br_13
port 30 nsew
rlabel metal1 s 7408 629 7408 629 4 br_10
port 24 nsew
rlabel metal1 s 18016 629 18016 629 4 bl_27
port 57 nsew
rlabel metal1 s 11152 629 11152 629 4 br_16
port 36 nsew
rlabel metal1 s 2576 629 2576 629 4 br_3
port 10 nsew
rlabel metal1 s 4912 629 4912 629 4 br_6
port 16 nsew
rlabel metal1 s 80 629 80 629 4 rbl_br
port 2 nsew
rlabel metal1 s 20048 629 20048 629 4 br_31
port 66 nsew
rlabel metal1 s 14272 629 14272 629 4 bl_21
port 45 nsew
rlabel metal1 s 3200 629 3200 629 4 bl_4
port 11 nsew
rlabel metal1 s 13648 629 13648 629 4 br_20
port 44 nsew
rlabel metal1 s 14896 629 14896 629 4 br_22
port 48 nsew
rlabel metal1 s 18640 629 18640 629 4 br_28
port 60 nsew
rlabel metal1 s 16304 629 16304 629 4 br_25
port 54 nsew
rlabel metal1 s 19264 629 19264 629 4 bl_29
port 61 nsew
rlabel metal1 s 15680 629 15680 629 4 bl_24
port 51 nsew
rlabel metal1 s 19888 629 19888 629 4 br_30
port 64 nsew
rlabel metal1 s 544 629 544 629 4 rbl_bl
port 1 nsew
rlabel metal1 s 13024 629 13024 629 4 bl_19
port 41 nsew
rlabel metal1 s 6160 629 6160 629 4 br_8
port 20 nsew
rlabel metal1 s 10528 629 10528 629 4 bl_15
port 33 nsew
rlabel metal1 s 6784 629 6784 629 4 bl_9
port 21 nsew
rlabel metal1 s 6320 629 6320 629 4 br_9
port 22 nsew
rlabel metal1 s 4288 629 4288 629 4 bl_5
port 13 nsew
rlabel metal1 s 16768 629 16768 629 4 bl_25
port 53 nsew
rlabel metal1 s 8032 629 8032 629 4 bl_11
port 25 nsew
rlabel metal1 s 6944 629 6944 629 4 bl_10
port 23 nsew
rlabel metal1 s 14432 629 14432 629 4 bl_22
port 47 nsew
rlabel metal1 s 10064 629 10064 629 4 br_15
port 34 nsew
rlabel metal1 s 3824 629 3824 629 4 br_5
port 14 nsew
rlabel metal1 s 12560 629 12560 629 4 br_19
port 42 nsew
rlabel metal1 s 9280 629 9280 629 4 bl_13
port 29 nsew
rlabel metal1 s 3664 629 3664 629 4 br_4
port 12 nsew
rlabel metal1 s 9904 629 9904 629 4 br_14
port 32 nsew
rlabel metal1 s 4448 629 4448 629 4 bl_6
port 15 nsew
rlabel metal1 s 1168 629 1168 629 4 br_0
port 4 nsew
rlabel metal1 s 16144 629 16144 629 4 br_24
port 52 nsew
rlabel metal1 s 17552 629 17552 629 4 br_27
port 58 nsew
rlabel metal1 s 2416 629 2416 629 4 br_2
port 8 nsew
rlabel metal1 s 18176 629 18176 629 4 bl_28
port 59 nsew
rlabel metal1 s 5072 629 5072 629 4 br_7
port 18 nsew
rlabel metal1 s 18800 629 18800 629 4 br_29
port 62 nsew
rlabel metal1 s 704 629 704 629 4 bl_0
port 3 nsew
rlabel metal1 s 9440 629 9440 629 4 bl_14
port 31 nsew
rlabel metal1 s 5696 629 5696 629 4 bl_8
port 19 nsew
rlabel metal1 s 26128 629 26128 629 4 br_40
port 84 nsew
rlabel metal1 s 38144 629 38144 629 4 bl_60
port 123 nsew
rlabel metal1 s 38608 629 38608 629 4 br_60
port 124 nsew
rlabel metal1 s 31904 629 31904 629 4 bl_50
port 103 nsew
rlabel metal1 s 39232 629 39232 629 4 bl_61
port 125 nsew
rlabel metal1 s 39856 629 39856 629 4 br_62
port 128 nsew
rlabel metal1 s 26288 629 26288 629 4 br_41
port 86 nsew
rlabel metal1 s 27536 629 27536 629 4 br_43
port 90 nsew
rlabel metal1 s 29248 629 29248 629 4 bl_45
port 93 nsew
rlabel metal1 s 24256 629 24256 629 4 bl_37
port 77 nsew
rlabel metal1 s 23792 629 23792 629 4 br_37
port 78 nsew
rlabel metal1 s 37984 629 37984 629 4 bl_59
port 121 nsew
rlabel metal1 s 36272 629 36272 629 4 br_57
port 118 nsew
rlabel metal1 s 28624 629 28624 629 4 br_44
port 92 nsew
rlabel metal1 s 22544 629 22544 629 4 br_35
port 74 nsew
rlabel metal1 s 34400 629 34400 629 4 bl_54
port 111 nsew
rlabel metal1 s 33616 629 33616 629 4 br_52
port 108 nsew
rlabel metal1 s 34240 629 34240 629 4 bl_53
port 109 nsew
rlabel metal1 s 34864 629 34864 629 4 br_54
port 112 nsew
rlabel metal1 s 33776 629 33776 629 4 br_53
port 110 nsew
rlabel metal1 s 24416 629 24416 629 4 bl_38
port 79 nsew
rlabel metal1 s 20672 629 20672 629 4 bl_32
port 67 nsew
rlabel metal1 s 35024 629 35024 629 4 br_55
port 114 nsew
rlabel metal1 s 37520 629 37520 629 4 br_59
port 122 nsew
rlabel metal1 s 29408 629 29408 629 4 bl_46
port 95 nsew
rlabel metal1 s 33152 629 33152 629 4 bl_52
port 107 nsew
rlabel metal1 s 28160 629 28160 629 4 bl_44
port 91 nsew
rlabel metal1 s 37360 629 37360 629 4 br_58
port 120 nsew
rlabel metal1 s 35488 629 35488 629 4 bl_55
port 113 nsew
rlabel metal1 s 35648 629 35648 629 4 bl_56
port 115 nsew
rlabel metal1 s 31744 629 31744 629 4 bl_49
port 101 nsew
rlabel metal1 s 28784 629 28784 629 4 br_45
port 94 nsew
rlabel metal1 s 23168 629 23168 629 4 bl_36
port 75 nsew
rlabel metal1 s 24880 629 24880 629 4 br_38
port 80 nsew
rlabel metal1 s 27376 629 27376 629 4 br_42
port 88 nsew
rlabel metal1 s 21136 629 21136 629 4 br_32
port 68 nsew
rlabel metal1 s 23008 629 23008 629 4 bl_35
port 73 nsew
rlabel metal1 s 31280 629 31280 629 4 br_49
port 102 nsew
rlabel metal1 s 40016 629 40016 629 4 br_63
port 130 nsew
rlabel metal1 s 29872 629 29872 629 4 br_46
port 96 nsew
rlabel metal1 s 20512 629 20512 629 4 bl_31
port 65 nsew
rlabel metal1 s 30032 629 30032 629 4 br_47
port 98 nsew
rlabel metal1 s 25664 629 25664 629 4 bl_40
port 83 nsew
rlabel metal1 s 30496 629 30496 629 4 bl_47
port 97 nsew
rlabel metal1 s 21760 629 21760 629 4 bl_33
port 69 nsew
rlabel metal1 s 22384 629 22384 629 4 br_34
port 72 nsew
rlabel metal1 s 39392 629 39392 629 4 bl_62
port 127 nsew
rlabel metal1 s 28000 629 28000 629 4 bl_43
port 89 nsew
rlabel metal1 s 26912 629 26912 629 4 bl_42
port 87 nsew
rlabel metal1 s 40480 629 40480 629 4 bl_63
port 129 nsew
rlabel metal1 s 30656 629 30656 629 4 bl_48
port 99 nsew
rlabel metal1 s 26752 629 26752 629 4 bl_41
port 85 nsew
rlabel metal1 s 25504 629 25504 629 4 bl_39
port 81 nsew
rlabel metal1 s 38768 629 38768 629 4 br_61
port 126 nsew
rlabel metal1 s 21296 629 21296 629 4 br_33
port 70 nsew
rlabel metal1 s 36896 629 36896 629 4 bl_58
port 119 nsew
rlabel metal1 s 25040 629 25040 629 4 br_39
port 82 nsew
rlabel metal1 s 23632 629 23632 629 4 br_36
port 76 nsew
rlabel metal1 s 32992 629 32992 629 4 bl_51
port 105 nsew
rlabel metal1 s 31120 629 31120 629 4 br_48
port 100 nsew
rlabel metal1 s 36736 629 36736 629 4 bl_57
port 117 nsew
rlabel metal1 s 21920 629 21920 629 4 bl_34
port 71 nsew
rlabel metal1 s 32368 629 32368 629 4 br_50
port 104 nsew
rlabel metal1 s 36112 629 36112 629 4 br_56
port 116 nsew
rlabel metal1 s 32528 629 32528 629 4 br_51
port 106 nsew
rlabel metal2 s 10608 9115 10608 9115 4 bank_wmask_1
port 73 nsew
rlabel metal2 s 624 9115 624 9115 4 bank_wmask_0
port 72 nsew
rlabel metal2 s 30576 9115 30576 9115 4 bank_wmask_3
port 75 nsew
rlabel metal2 s 20592 9115 20592 9115 4 bank_wmask_2
port 74 nsew
rlabel metal3 s 34697 7204 34697 7204 4 gnd
port 77 nsew
rlabel metal3 s 39574 7406 39574 7406 4 gnd
port 77 nsew
rlabel metal3 s 35945 7204 35945 7204 4 gnd
port 77 nsew
rlabel metal3 s 30949 9385 30949 9385 4 gnd
port 77 nsew
rlabel metal3 s 34582 7406 34582 7406 4 gnd
port 77 nsew
rlabel metal3 s 32086 7406 32086 7406 4 gnd
port 77 nsew
rlabel metal3 s 39689 7204 39689 7204 4 gnd
port 77 nsew
rlabel metal3 s 33334 7406 33334 7406 4 gnd
port 77 nsew
rlabel metal3 s 35830 7406 35830 7406 4 gnd
port 77 nsew
rlabel metal3 s 30838 7406 30838 7406 4 gnd
port 77 nsew
rlabel metal3 s 33449 7204 33449 7204 4 gnd
port 77 nsew
rlabel metal3 s 37193 7204 37193 7204 4 gnd
port 77 nsew
rlabel metal3 s 37078 7406 37078 7406 4 gnd
port 77 nsew
rlabel metal3 s 32201 7204 32201 7204 4 gnd
port 77 nsew
rlabel metal3 s 38326 7406 38326 7406 4 gnd
port 77 nsew
rlabel metal3 s 38441 7204 38441 7204 4 gnd
port 77 nsew
rlabel metal3 s 30953 7204 30953 7204 4 gnd
port 77 nsew
rlabel metal3 s 33348 7822 33348 7822 4 vdd
port 76 nsew
rlabel metal3 s 30949 8265 30949 8265 4 vdd
port 76 nsew
rlabel metal3 s 39588 7822 39588 7822 4 vdd
port 76 nsew
rlabel metal3 s 37092 7822 37092 7822 4 vdd
port 76 nsew
rlabel metal3 s 35844 7822 35844 7822 4 vdd
port 76 nsew
rlabel metal3 s 38340 7822 38340 7822 4 vdd
port 76 nsew
rlabel metal3 s 30852 7822 30852 7822 4 vdd
port 76 nsew
rlabel metal3 s 34596 7822 34596 7822 4 vdd
port 76 nsew
rlabel metal3 s 32100 7822 32100 7822 4 vdd
port 76 nsew
rlabel metal3 s 35949 5642 35949 5642 4 gnd
port 77 nsew
rlabel metal3 s 35835 6435 35835 6435 4 gnd
port 77 nsew
rlabel metal3 s 39693 5642 39693 5642 4 gnd
port 77 nsew
rlabel metal3 s 37072 6872 37072 6872 4 vdd
port 76 nsew
rlabel metal3 s 38445 5642 38445 5642 4 gnd
port 77 nsew
rlabel metal3 s 38331 6435 38331 6435 4 gnd
port 77 nsew
rlabel metal3 s 32205 5642 32205 5642 4 gnd
port 77 nsew
rlabel metal3 s 33453 5642 33453 5642 4 gnd
port 77 nsew
rlabel metal3 s 30957 5642 30957 5642 4 gnd
port 77 nsew
rlabel metal3 s 32205 5320 32205 5320 4 vdd
port 76 nsew
rlabel metal3 s 37197 5642 37197 5642 4 gnd
port 77 nsew
rlabel metal3 s 30843 6435 30843 6435 4 gnd
port 77 nsew
rlabel metal3 s 33339 6435 33339 6435 4 gnd
port 77 nsew
rlabel metal3 s 38445 5320 38445 5320 4 vdd
port 76 nsew
rlabel metal3 s 35824 6872 35824 6872 4 vdd
port 76 nsew
rlabel metal3 s 33328 6872 33328 6872 4 vdd
port 76 nsew
rlabel metal3 s 38320 6872 38320 6872 4 vdd
port 76 nsew
rlabel metal3 s 37197 5320 37197 5320 4 vdd
port 76 nsew
rlabel metal3 s 33453 5320 33453 5320 4 vdd
port 76 nsew
rlabel metal3 s 34587 6435 34587 6435 4 gnd
port 77 nsew
rlabel metal3 s 30957 5320 30957 5320 4 vdd
port 76 nsew
rlabel metal3 s 35949 5320 35949 5320 4 vdd
port 76 nsew
rlabel metal3 s 34576 6872 34576 6872 4 vdd
port 76 nsew
rlabel metal3 s 34701 5642 34701 5642 4 gnd
port 77 nsew
rlabel metal3 s 39579 6435 39579 6435 4 gnd
port 77 nsew
rlabel metal3 s 39693 5320 39693 5320 4 vdd
port 76 nsew
rlabel metal3 s 34701 5320 34701 5320 4 vdd
port 76 nsew
rlabel metal3 s 32091 6435 32091 6435 4 gnd
port 77 nsew
rlabel metal3 s 39568 6872 39568 6872 4 vdd
port 76 nsew
rlabel metal3 s 32080 6872 32080 6872 4 vdd
port 76 nsew
rlabel metal3 s 30832 6872 30832 6872 4 vdd
port 76 nsew
rlabel metal3 s 37083 6435 37083 6435 4 gnd
port 77 nsew
rlabel metal3 s 22096 6872 22096 6872 4 vdd
port 76 nsew
rlabel metal3 s 22221 5642 22221 5642 4 gnd
port 77 nsew
rlabel metal3 s 24592 6872 24592 6872 4 vdd
port 76 nsew
rlabel metal3 s 22221 5320 22221 5320 4 vdd
port 76 nsew
rlabel metal3 s 29595 6435 29595 6435 4 gnd
port 77 nsew
rlabel metal3 s 27213 5642 27213 5642 4 gnd
port 77 nsew
rlabel metal3 s 27099 6435 27099 6435 4 gnd
port 77 nsew
rlabel metal3 s 25965 5642 25965 5642 4 gnd
port 77 nsew
rlabel metal3 s 23355 6435 23355 6435 4 gnd
port 77 nsew
rlabel metal3 s 20848 6872 20848 6872 4 vdd
port 76 nsew
rlabel metal3 s 28461 5320 28461 5320 4 vdd
port 76 nsew
rlabel metal3 s 24717 5642 24717 5642 4 gnd
port 77 nsew
rlabel metal3 s 29709 5642 29709 5642 4 gnd
port 77 nsew
rlabel metal3 s 25840 6872 25840 6872 4 vdd
port 76 nsew
rlabel metal3 s 23469 5320 23469 5320 4 vdd
port 76 nsew
rlabel metal3 s 28461 5642 28461 5642 4 gnd
port 77 nsew
rlabel metal3 s 22107 6435 22107 6435 4 gnd
port 77 nsew
rlabel metal3 s 24603 6435 24603 6435 4 gnd
port 77 nsew
rlabel metal3 s 27088 6872 27088 6872 4 vdd
port 76 nsew
rlabel metal3 s 23469 5642 23469 5642 4 gnd
port 77 nsew
rlabel metal3 s 27213 5320 27213 5320 4 vdd
port 76 nsew
rlabel metal3 s 23344 6872 23344 6872 4 vdd
port 76 nsew
rlabel metal3 s 20973 5642 20973 5642 4 gnd
port 77 nsew
rlabel metal3 s 20973 5320 20973 5320 4 vdd
port 76 nsew
rlabel metal3 s 29709 5320 29709 5320 4 vdd
port 76 nsew
rlabel metal3 s 20859 6435 20859 6435 4 gnd
port 77 nsew
rlabel metal3 s 28336 6872 28336 6872 4 vdd
port 76 nsew
rlabel metal3 s 20854 7406 20854 7406 4 gnd
port 77 nsew
rlabel metal3 s 29705 7204 29705 7204 4 gnd
port 77 nsew
rlabel metal3 s 22217 7204 22217 7204 4 gnd
port 77 nsew
rlabel metal3 s 20969 7204 20969 7204 4 gnd
port 77 nsew
rlabel metal3 s 27094 7406 27094 7406 4 gnd
port 77 nsew
rlabel metal3 s 27209 7204 27209 7204 4 gnd
port 77 nsew
rlabel metal3 s 28342 7406 28342 7406 4 gnd
port 77 nsew
rlabel metal3 s 25846 7406 25846 7406 4 gnd
port 77 nsew
rlabel metal3 s 28457 7204 28457 7204 4 gnd
port 77 nsew
rlabel metal3 s 24713 7204 24713 7204 4 gnd
port 77 nsew
rlabel metal3 s 29590 7406 29590 7406 4 gnd
port 77 nsew
rlabel metal3 s 25860 7822 25860 7822 4 vdd
port 76 nsew
rlabel metal3 s 25961 7204 25961 7204 4 gnd
port 77 nsew
rlabel metal3 s 22102 7406 22102 7406 4 gnd
port 77 nsew
rlabel metal3 s 20965 9385 20965 9385 4 gnd
port 77 nsew
rlabel metal3 s 23350 7406 23350 7406 4 gnd
port 77 nsew
rlabel metal3 s 23364 7822 23364 7822 4 vdd
port 76 nsew
rlabel metal3 s 20592 8867 20592 8867 4 w_en
port 71 nsew
rlabel metal3 s 22116 7822 22116 7822 4 vdd
port 76 nsew
rlabel metal3 s 29604 7822 29604 7822 4 vdd
port 76 nsew
rlabel metal3 s 24612 7822 24612 7822 4 vdd
port 76 nsew
rlabel metal3 s 23465 7204 23465 7204 4 gnd
port 77 nsew
rlabel metal3 s 20965 8265 20965 8265 4 vdd
port 76 nsew
rlabel metal3 s 27108 7822 27108 7822 4 vdd
port 76 nsew
rlabel metal3 s 28356 7822 28356 7822 4 vdd
port 76 nsew
rlabel metal3 s 20868 7822 20868 7822 4 vdd
port 76 nsew
rlabel metal3 s 24598 7406 24598 7406 4 gnd
port 77 nsew
rlabel metal3 s 25851 6435 25851 6435 4 gnd
port 77 nsew
rlabel metal3 s 25965 5320 25965 5320 4 vdd
port 76 nsew
rlabel metal3 s 24717 5320 24717 5320 4 vdd
port 76 nsew
rlabel metal3 s 28347 6435 28347 6435 4 gnd
port 77 nsew
rlabel metal3 s 29584 6872 29584 6872 4 vdd
port 76 nsew
rlabel metal3 s 28704 1935 28704 1935 4 gnd
port 77 nsew
rlabel metal3 s 23539 3708 23539 3708 4 gnd
port 77 nsew
rlabel metal3 s 26208 1935 26208 1935 4 gnd
port 77 nsew
rlabel metal3 s 23712 1935 23712 1935 4 gnd
port 77 nsew
rlabel metal3 s 23457 4482 23457 4482 4 vdd
port 76 nsew
rlabel metal3 s 29779 3708 29779 3708 4 gnd
port 77 nsew
rlabel metal3 s 22464 1935 22464 1935 4 gnd
port 77 nsew
rlabel metal3 s 24787 3708 24787 3708 4 gnd
port 77 nsew
rlabel metal3 s 22209 4482 22209 4482 4 vdd
port 76 nsew
rlabel metal3 s 28449 4482 28449 4482 4 vdd
port 76 nsew
rlabel metal3 s 27283 3708 27283 3708 4 gnd
port 77 nsew
rlabel metal3 s 29697 4482 29697 4482 4 vdd
port 76 nsew
rlabel metal3 s 25953 4482 25953 4482 4 vdd
port 76 nsew
rlabel metal3 s 29952 1935 29952 1935 4 gnd
port 77 nsew
rlabel metal3 s 24960 1935 24960 1935 4 gnd
port 77 nsew
rlabel metal3 s 20592 3556 20592 3556 4 s_en
port 69 nsew
rlabel metal3 s 20592 2840 20592 2840 4 sel_0
port 67 nsew
rlabel metal3 s 22291 3708 22291 3708 4 gnd
port 77 nsew
rlabel metal3 s 27456 1935 27456 1935 4 gnd
port 77 nsew
rlabel metal3 s 27201 4482 27201 4482 4 vdd
port 76 nsew
rlabel metal3 s 21216 1935 21216 1935 4 gnd
port 77 nsew
rlabel metal3 s 28531 3708 28531 3708 4 gnd
port 77 nsew
rlabel metal3 s 20961 4482 20961 4482 4 vdd
port 76 nsew
rlabel metal3 s 26035 3708 26035 3708 4 gnd
port 77 nsew
rlabel metal3 s 24705 4482 24705 4482 4 vdd
port 76 nsew
rlabel metal3 s 21043 3708 21043 3708 4 gnd
port 77 nsew
rlabel metal3 s 20592 2716 20592 2716 4 sel_1
port 68 nsew
rlabel metal3 s 39763 3708 39763 3708 4 gnd
port 77 nsew
rlabel metal3 s 37267 3708 37267 3708 4 gnd
port 77 nsew
rlabel metal3 s 39936 1935 39936 1935 4 gnd
port 77 nsew
rlabel metal3 s 37185 4482 37185 4482 4 vdd
port 76 nsew
rlabel metal3 s 35937 4482 35937 4482 4 vdd
port 76 nsew
rlabel metal3 s 33696 1935 33696 1935 4 gnd
port 77 nsew
rlabel metal3 s 31200 1935 31200 1935 4 gnd
port 77 nsew
rlabel metal3 s 32193 4482 32193 4482 4 vdd
port 76 nsew
rlabel metal3 s 32448 1935 32448 1935 4 gnd
port 77 nsew
rlabel metal3 s 38515 3708 38515 3708 4 gnd
port 77 nsew
rlabel metal3 s 37440 1935 37440 1935 4 gnd
port 77 nsew
rlabel metal3 s 33441 4482 33441 4482 4 vdd
port 76 nsew
rlabel metal3 s 31027 3708 31027 3708 4 gnd
port 77 nsew
rlabel metal3 s 36019 3708 36019 3708 4 gnd
port 77 nsew
rlabel metal3 s 38433 4482 38433 4482 4 vdd
port 76 nsew
rlabel metal3 s 39681 4482 39681 4482 4 vdd
port 76 nsew
rlabel metal3 s 34689 4482 34689 4482 4 vdd
port 76 nsew
rlabel metal3 s 32275 3708 32275 3708 4 gnd
port 77 nsew
rlabel metal3 s 34944 1935 34944 1935 4 gnd
port 77 nsew
rlabel metal3 s 30945 4482 30945 4482 4 vdd
port 76 nsew
rlabel metal3 s 34771 3708 34771 3708 4 gnd
port 77 nsew
rlabel metal3 s 36192 1935 36192 1935 4 gnd
port 77 nsew
rlabel metal3 s 38688 1935 38688 1935 4 gnd
port 77 nsew
rlabel metal3 s 33523 3708 33523 3708 4 gnd
port 77 nsew
rlabel metal3 s 14608 6872 14608 6872 4 vdd
port 76 nsew
rlabel metal3 s 18477 5320 18477 5320 4 vdd
port 76 nsew
rlabel metal3 s 17115 6435 17115 6435 4 gnd
port 77 nsew
rlabel metal3 s 10875 6435 10875 6435 4 gnd
port 77 nsew
rlabel metal3 s 17229 5320 17229 5320 4 vdd
port 76 nsew
rlabel metal3 s 15981 5642 15981 5642 4 gnd
port 77 nsew
rlabel metal3 s 17104 6872 17104 6872 4 vdd
port 76 nsew
rlabel metal3 s 14733 5642 14733 5642 4 gnd
port 77 nsew
rlabel metal3 s 10989 5320 10989 5320 4 vdd
port 76 nsew
rlabel metal3 s 17229 5642 17229 5642 4 gnd
port 77 nsew
rlabel metal3 s 13485 5642 13485 5642 4 gnd
port 77 nsew
rlabel metal3 s 10864 6872 10864 6872 4 vdd
port 76 nsew
rlabel metal3 s 13360 6872 13360 6872 4 vdd
port 76 nsew
rlabel metal3 s 12112 6872 12112 6872 4 vdd
port 76 nsew
rlabel metal3 s 18363 6435 18363 6435 4 gnd
port 77 nsew
rlabel metal3 s 13371 6435 13371 6435 4 gnd
port 77 nsew
rlabel metal3 s 12237 5642 12237 5642 4 gnd
port 77 nsew
rlabel metal3 s 19611 6435 19611 6435 4 gnd
port 77 nsew
rlabel metal3 s 18352 6872 18352 6872 4 vdd
port 76 nsew
rlabel metal3 s 12123 6435 12123 6435 4 gnd
port 77 nsew
rlabel metal3 s 19600 6872 19600 6872 4 vdd
port 76 nsew
rlabel metal3 s 19725 5320 19725 5320 4 vdd
port 76 nsew
rlabel metal3 s 14619 6435 14619 6435 4 gnd
port 77 nsew
rlabel metal3 s 15981 5320 15981 5320 4 vdd
port 76 nsew
rlabel metal3 s 15856 6872 15856 6872 4 vdd
port 76 nsew
rlabel metal3 s 15867 6435 15867 6435 4 gnd
port 77 nsew
rlabel metal3 s 13485 5320 13485 5320 4 vdd
port 76 nsew
rlabel metal3 s 18477 5642 18477 5642 4 gnd
port 77 nsew
rlabel metal3 s 14733 5320 14733 5320 4 vdd
port 76 nsew
rlabel metal3 s 12237 5320 12237 5320 4 vdd
port 76 nsew
rlabel metal3 s 10989 5642 10989 5642 4 gnd
port 77 nsew
rlabel metal3 s 19725 5642 19725 5642 4 gnd
port 77 nsew
rlabel metal3 s 14614 7406 14614 7406 4 gnd
port 77 nsew
rlabel metal3 s 12118 7406 12118 7406 4 gnd
port 77 nsew
rlabel metal3 s 15862 7406 15862 7406 4 gnd
port 77 nsew
rlabel metal3 s 19606 7406 19606 7406 4 gnd
port 77 nsew
rlabel metal3 s 13366 7406 13366 7406 4 gnd
port 77 nsew
rlabel metal3 s 10981 8265 10981 8265 4 vdd
port 76 nsew
rlabel metal3 s 12132 7822 12132 7822 4 vdd
port 76 nsew
rlabel metal3 s 12233 7204 12233 7204 4 gnd
port 77 nsew
rlabel metal3 s 17110 7406 17110 7406 4 gnd
port 77 nsew
rlabel metal3 s 18372 7822 18372 7822 4 vdd
port 76 nsew
rlabel metal3 s 18473 7204 18473 7204 4 gnd
port 77 nsew
rlabel metal3 s 14628 7822 14628 7822 4 vdd
port 76 nsew
rlabel metal3 s 10884 7822 10884 7822 4 vdd
port 76 nsew
rlabel metal3 s 15977 7204 15977 7204 4 gnd
port 77 nsew
rlabel metal3 s 19620 7822 19620 7822 4 vdd
port 76 nsew
rlabel metal3 s 10870 7406 10870 7406 4 gnd
port 77 nsew
rlabel metal3 s 10981 9385 10981 9385 4 gnd
port 77 nsew
rlabel metal3 s 17225 7204 17225 7204 4 gnd
port 77 nsew
rlabel metal3 s 10985 7204 10985 7204 4 gnd
port 77 nsew
rlabel metal3 s 18358 7406 18358 7406 4 gnd
port 77 nsew
rlabel metal3 s 19721 7204 19721 7204 4 gnd
port 77 nsew
rlabel metal3 s 17124 7822 17124 7822 4 vdd
port 76 nsew
rlabel metal3 s 13380 7822 13380 7822 4 vdd
port 76 nsew
rlabel metal3 s 15876 7822 15876 7822 4 vdd
port 76 nsew
rlabel metal3 s 14729 7204 14729 7204 4 gnd
port 77 nsew
rlabel metal3 s 13481 7204 13481 7204 4 gnd
port 77 nsew
rlabel metal3 s 8379 6435 8379 6435 4 gnd
port 77 nsew
rlabel metal3 s 9616 6872 9616 6872 4 vdd
port 76 nsew
rlabel metal3 s 4749 5320 4749 5320 4 vdd
port 76 nsew
rlabel metal3 s 8493 5642 8493 5642 4 gnd
port 77 nsew
rlabel metal3 s 891 6435 891 6435 4 gnd
port 77 nsew
rlabel metal3 s 7131 6435 7131 6435 4 gnd
port 77 nsew
rlabel metal3 s 4635 6435 4635 6435 4 gnd
port 77 nsew
rlabel metal3 s 4749 5642 4749 5642 4 gnd
port 77 nsew
rlabel metal3 s 3382 7406 3382 7406 4 gnd
port 77 nsew
rlabel metal3 s 2139 6435 2139 6435 4 gnd
port 77 nsew
rlabel metal3 s 3501 5642 3501 5642 4 gnd
port 77 nsew
rlabel metal3 s 8493 5320 8493 5320 4 vdd
port 76 nsew
rlabel metal3 s 9741 5642 9741 5642 4 gnd
port 77 nsew
rlabel metal3 s 2128 6872 2128 6872 4 vdd
port 76 nsew
rlabel metal3 s 9741 5320 9741 5320 4 vdd
port 76 nsew
rlabel metal3 s 7245 5642 7245 5642 4 gnd
port 77 nsew
rlabel metal3 s 880 6872 880 6872 4 vdd
port 76 nsew
rlabel metal3 s 2253 5642 2253 5642 4 gnd
port 77 nsew
rlabel metal3 s 5872 6872 5872 6872 4 vdd
port 76 nsew
rlabel metal3 s 3376 6872 3376 6872 4 vdd
port 76 nsew
rlabel metal3 s 5997 5320 5997 5320 4 vdd
port 76 nsew
rlabel metal3 s 2253 5320 2253 5320 4 vdd
port 76 nsew
rlabel metal3 s 8368 6872 8368 6872 4 vdd
port 76 nsew
rlabel metal3 s 7120 6872 7120 6872 4 vdd
port 76 nsew
rlabel metal3 s 1005 5320 1005 5320 4 vdd
port 76 nsew
rlabel metal3 s 5997 5642 5997 5642 4 gnd
port 77 nsew
rlabel metal3 s 9627 6435 9627 6435 4 gnd
port 77 nsew
rlabel metal3 s 3387 6435 3387 6435 4 gnd
port 77 nsew
rlabel metal3 s 5883 6435 5883 6435 4 gnd
port 77 nsew
rlabel metal3 s 3501 5320 3501 5320 4 vdd
port 76 nsew
rlabel metal3 s 7245 5320 7245 5320 4 vdd
port 76 nsew
rlabel metal3 s 4624 6872 4624 6872 4 vdd
port 76 nsew
rlabel metal3 s 1005 5642 1005 5642 4 gnd
port 77 nsew
rlabel metal3 s 9636 7822 9636 7822 4 vdd
port 76 nsew
rlabel metal3 s 7140 7822 7140 7822 4 vdd
port 76 nsew
rlabel metal3 s 886 7406 886 7406 4 gnd
port 77 nsew
rlabel metal3 s 1001 7204 1001 7204 4 gnd
port 77 nsew
rlabel metal3 s 5993 7204 5993 7204 4 gnd
port 77 nsew
rlabel metal3 s 7241 7204 7241 7204 4 gnd
port 77 nsew
rlabel metal3 s 997 9385 997 9385 4 gnd
port 77 nsew
rlabel metal3 s 3396 7822 3396 7822 4 vdd
port 76 nsew
rlabel metal3 s 997 8265 997 8265 4 vdd
port 76 nsew
rlabel metal3 s 4630 7406 4630 7406 4 gnd
port 77 nsew
rlabel metal3 s 4745 7204 4745 7204 4 gnd
port 77 nsew
rlabel metal3 s 8489 7204 8489 7204 4 gnd
port 77 nsew
rlabel metal3 s 5892 7822 5892 7822 4 vdd
port 76 nsew
rlabel metal3 s 2134 7406 2134 7406 4 gnd
port 77 nsew
rlabel metal3 s 7126 7406 7126 7406 4 gnd
port 77 nsew
rlabel metal3 s 8374 7406 8374 7406 4 gnd
port 77 nsew
rlabel metal3 s 5878 7406 5878 7406 4 gnd
port 77 nsew
rlabel metal3 s 4644 7822 4644 7822 4 vdd
port 76 nsew
rlabel metal3 s 8388 7822 8388 7822 4 vdd
port 76 nsew
rlabel metal3 s 9737 7204 9737 7204 4 gnd
port 77 nsew
rlabel metal3 s 900 7822 900 7822 4 vdd
port 76 nsew
rlabel metal3 s 9622 7406 9622 7406 4 gnd
port 77 nsew
rlabel metal3 s 3497 7204 3497 7204 4 gnd
port 77 nsew
rlabel metal3 s 2249 7204 2249 7204 4 gnd
port 77 nsew
rlabel metal3 s 2148 7822 2148 7822 4 vdd
port 76 nsew
rlabel metal3 s 4819 3708 4819 3708 4 gnd
port 77 nsew
rlabel metal3 s 8736 1935 8736 1935 4 gnd
port 77 nsew
rlabel metal3 s 6240 1935 6240 1935 4 gnd
port 77 nsew
rlabel metal3 s 7315 3708 7315 3708 4 gnd
port 77 nsew
rlabel metal3 s 1248 1935 1248 1935 4 gnd
port 77 nsew
rlabel metal3 s 3489 4482 3489 4482 4 vdd
port 76 nsew
rlabel metal3 s 4992 1935 4992 1935 4 gnd
port 77 nsew
rlabel metal3 s 9984 1935 9984 1935 4 gnd
port 77 nsew
rlabel metal3 s 2496 1935 2496 1935 4 gnd
port 77 nsew
rlabel metal3 s 2323 3708 2323 3708 4 gnd
port 77 nsew
rlabel metal3 s 2241 4482 2241 4482 4 vdd
port 76 nsew
rlabel metal3 s 9729 4482 9729 4482 4 vdd
port 76 nsew
rlabel metal3 s 8563 3708 8563 3708 4 gnd
port 77 nsew
rlabel metal3 s 1075 3708 1075 3708 4 gnd
port 77 nsew
rlabel metal3 s 7488 1935 7488 1935 4 gnd
port 77 nsew
rlabel metal3 s 7233 4482 7233 4482 4 vdd
port 76 nsew
rlabel metal3 s 3744 1935 3744 1935 4 gnd
port 77 nsew
rlabel metal3 s 3571 3708 3571 3708 4 gnd
port 77 nsew
rlabel metal3 s 4737 4482 4737 4482 4 vdd
port 76 nsew
rlabel metal3 s 993 4482 993 4482 4 vdd
port 76 nsew
rlabel metal3 s 8481 4482 8481 4482 4 vdd
port 76 nsew
rlabel metal3 s 6067 3708 6067 3708 4 gnd
port 77 nsew
rlabel metal3 s 9811 3708 9811 3708 4 gnd
port 77 nsew
rlabel metal3 s 5985 4482 5985 4482 4 vdd
port 76 nsew
rlabel metal3 s 18465 4482 18465 4482 4 vdd
port 76 nsew
rlabel metal3 s 17299 3708 17299 3708 4 gnd
port 77 nsew
rlabel metal3 s 13473 4482 13473 4482 4 vdd
port 76 nsew
rlabel metal3 s 13728 1935 13728 1935 4 gnd
port 77 nsew
rlabel metal3 s 14721 4482 14721 4482 4 vdd
port 76 nsew
rlabel metal3 s 14976 1935 14976 1935 4 gnd
port 77 nsew
rlabel metal3 s 16224 1935 16224 1935 4 gnd
port 77 nsew
rlabel metal3 s 18547 3708 18547 3708 4 gnd
port 77 nsew
rlabel metal3 s 16051 3708 16051 3708 4 gnd
port 77 nsew
rlabel metal3 s 11232 1935 11232 1935 4 gnd
port 77 nsew
rlabel metal3 s 14803 3708 14803 3708 4 gnd
port 77 nsew
rlabel metal3 s 11059 3708 11059 3708 4 gnd
port 77 nsew
rlabel metal3 s 10977 4482 10977 4482 4 vdd
port 76 nsew
rlabel metal3 s 18720 1935 18720 1935 4 gnd
port 77 nsew
rlabel metal3 s 19713 4482 19713 4482 4 vdd
port 76 nsew
rlabel metal3 s 19795 3708 19795 3708 4 gnd
port 77 nsew
rlabel metal3 s 17217 4482 17217 4482 4 vdd
port 76 nsew
rlabel metal3 s 12480 1935 12480 1935 4 gnd
port 77 nsew
rlabel metal3 s 15969 4482 15969 4482 4 vdd
port 76 nsew
rlabel metal3 s 12225 4482 12225 4482 4 vdd
port 76 nsew
rlabel metal3 s 19968 1935 19968 1935 4 gnd
port 77 nsew
rlabel metal3 s 20280 981 20280 981 4 p_en_bar
port 70 nsew
rlabel metal3 s 13555 3708 13555 3708 4 gnd
port 77 nsew
rlabel metal3 s 17472 1935 17472 1935 4 gnd
port 77 nsew
rlabel metal3 s 12307 3708 12307 3708 4 gnd
port 77 nsew
rlabel metal3 s 2927 362 2927 362 4 vdd
port 76 nsew
rlabel metal3 s 17041 362 17041 362 4 vdd
port 76 nsew
rlabel metal3 s 9553 362 9553 362 4 vdd
port 76 nsew
rlabel metal3 s 7919 362 7919 362 4 vdd
port 76 nsew
rlabel metal3 s 1679 362 1679 362 4 vdd
port 76 nsew
rlabel metal3 s 15407 362 15407 362 4 vdd
port 76 nsew
rlabel metal3 s 10801 362 10801 362 4 vdd
port 76 nsew
rlabel metal3 s 15793 362 15793 362 4 vdd
port 76 nsew
rlabel metal3 s 4175 362 4175 362 4 vdd
port 76 nsew
rlabel metal3 s 11663 362 11663 362 4 vdd
port 76 nsew
rlabel metal3 s 6671 362 6671 362 4 vdd
port 76 nsew
rlabel metal3 s 14545 362 14545 362 4 vdd
port 76 nsew
rlabel metal3 s 9167 362 9167 362 4 vdd
port 76 nsew
rlabel metal3 s 5423 362 5423 362 4 vdd
port 76 nsew
rlabel metal3 s 7057 362 7057 362 4 vdd
port 76 nsew
rlabel metal3 s 13297 362 13297 362 4 vdd
port 76 nsew
rlabel metal3 s 19537 362 19537 362 4 vdd
port 76 nsew
rlabel metal3 s 4561 362 4561 362 4 vdd
port 76 nsew
rlabel metal3 s 17903 362 17903 362 4 vdd
port 76 nsew
rlabel metal3 s 817 362 817 362 4 vdd
port 76 nsew
rlabel metal3 s 18289 362 18289 362 4 vdd
port 76 nsew
rlabel metal3 s 12049 362 12049 362 4 vdd
port 76 nsew
rlabel metal3 s 12911 362 12911 362 4 vdd
port 76 nsew
rlabel metal3 s 14159 362 14159 362 4 vdd
port 76 nsew
rlabel metal3 s 20399 362 20399 362 4 vdd
port 76 nsew
rlabel metal3 s 8305 362 8305 362 4 vdd
port 76 nsew
rlabel metal3 s 16655 362 16655 362 4 vdd
port 76 nsew
rlabel metal3 s 2065 362 2065 362 4 vdd
port 76 nsew
rlabel metal3 s 19151 362 19151 362 4 vdd
port 76 nsew
rlabel metal3 s 431 362 431 362 4 vdd
port 76 nsew
rlabel metal3 s 5809 362 5809 362 4 vdd
port 76 nsew
rlabel metal3 s 10415 362 10415 362 4 vdd
port 76 nsew
rlabel metal3 s 3313 362 3313 362 4 vdd
port 76 nsew
rlabel metal3 s 30769 362 30769 362 4 vdd
port 76 nsew
rlabel metal3 s 26639 362 26639 362 4 vdd
port 76 nsew
rlabel metal3 s 20785 362 20785 362 4 vdd
port 76 nsew
rlabel metal3 s 24143 362 24143 362 4 vdd
port 76 nsew
rlabel metal3 s 30383 362 30383 362 4 vdd
port 76 nsew
rlabel metal3 s 25391 362 25391 362 4 vdd
port 76 nsew
rlabel metal3 s 29521 362 29521 362 4 vdd
port 76 nsew
rlabel metal3 s 35761 362 35761 362 4 vdd
port 76 nsew
rlabel metal3 s 32879 362 32879 362 4 vdd
port 76 nsew
rlabel metal3 s 40367 362 40367 362 4 vdd
port 76 nsew
rlabel metal3 s 33265 362 33265 362 4 vdd
port 76 nsew
rlabel metal3 s 27025 362 27025 362 4 vdd
port 76 nsew
rlabel metal3 s 27887 362 27887 362 4 vdd
port 76 nsew
rlabel metal3 s 35375 362 35375 362 4 vdd
port 76 nsew
rlabel metal3 s 21647 362 21647 362 4 vdd
port 76 nsew
rlabel metal3 s 37871 362 37871 362 4 vdd
port 76 nsew
rlabel metal3 s 31631 362 31631 362 4 vdd
port 76 nsew
rlabel metal3 s 32017 362 32017 362 4 vdd
port 76 nsew
rlabel metal3 s 34513 362 34513 362 4 vdd
port 76 nsew
rlabel metal3 s 22895 362 22895 362 4 vdd
port 76 nsew
rlabel metal3 s 29135 362 29135 362 4 vdd
port 76 nsew
rlabel metal3 s 28273 362 28273 362 4 vdd
port 76 nsew
rlabel metal3 s 34127 362 34127 362 4 vdd
port 76 nsew
rlabel metal3 s 39505 362 39505 362 4 vdd
port 76 nsew
rlabel metal3 s 25777 362 25777 362 4 vdd
port 76 nsew
rlabel metal3 s 23281 362 23281 362 4 vdd
port 76 nsew
rlabel metal3 s 39119 362 39119 362 4 vdd
port 76 nsew
rlabel metal3 s 24529 362 24529 362 4 vdd
port 76 nsew
rlabel metal3 s 38257 362 38257 362 4 vdd
port 76 nsew
rlabel metal3 s 22033 362 22033 362 4 vdd
port 76 nsew
rlabel metal3 s 37009 362 37009 362 4 vdd
port 76 nsew
rlabel metal3 s 36623 362 36623 362 4 vdd
port 76 nsew
<< properties >>
string FIXED_BBOX 0 0 40560 9385
string GDS_END 4736336
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4578914
<< end >>
