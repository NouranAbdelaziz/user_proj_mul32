/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/parasitics/sky130_fd_pr__model__parasitic__rf_diode_ps2nw.model.spice