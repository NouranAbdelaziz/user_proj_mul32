magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
rect 222 0 258 52140
rect 294 0 330 52140
rect 366 51429 402 51770
rect 366 50639 402 51271
rect 366 49849 402 50481
rect 366 49059 402 49691
rect 366 48269 402 48901
rect 366 47479 402 48111
rect 366 46689 402 47321
rect 366 45899 402 46531
rect 366 45109 402 45741
rect 366 44319 402 44951
rect 366 43529 402 44161
rect 366 42739 402 43371
rect 366 41949 402 42581
rect 366 41159 402 41791
rect 366 40369 402 41001
rect 366 39579 402 40211
rect 366 38789 402 39421
rect 366 37999 402 38631
rect 366 37209 402 37841
rect 366 36419 402 37051
rect 366 35629 402 36261
rect 366 34839 402 35471
rect 366 34049 402 34681
rect 366 33259 402 33891
rect 366 32469 402 33101
rect 366 31679 402 32311
rect 366 30889 402 31521
rect 366 30099 402 30731
rect 366 29309 402 29941
rect 366 28519 402 29151
rect 366 27729 402 28361
rect 366 26939 402 27571
rect 366 26149 402 26781
rect 366 25359 402 25991
rect 366 24569 402 25201
rect 366 23779 402 24411
rect 366 22989 402 23621
rect 366 22199 402 22831
rect 366 21409 402 22041
rect 366 20619 402 21251
rect 366 19829 402 20461
rect 366 19039 402 19671
rect 366 18249 402 18881
rect 366 17459 402 18091
rect 366 16669 402 17301
rect 366 15879 402 16511
rect 366 15089 402 15721
rect 366 14299 402 14931
rect 366 13509 402 14141
rect 366 12719 402 13351
rect 366 11929 402 12561
rect 366 11139 402 11771
rect 366 10349 402 10981
rect 366 9559 402 10191
rect 366 8769 402 9401
rect 366 7979 402 8611
rect 366 7189 402 7821
rect 366 6399 402 7031
rect 366 5609 402 6241
rect 366 4819 402 5451
rect 366 4029 402 4661
rect 366 3239 402 3871
rect 366 2449 402 3081
rect 366 1659 402 2291
rect 366 869 402 1501
rect 366 370 402 711
rect 438 0 474 52140
rect 510 0 546 52140
<< metal2 >>
rect 284 51939 340 51948
rect 284 51874 340 51883
rect 0 51673 624 51721
rect 330 51549 438 51625
rect 0 51453 624 51501
rect 330 51295 438 51405
rect 0 51199 624 51247
rect 330 51075 438 51151
rect 0 50979 624 51027
rect 0 50883 624 50931
rect 330 50759 438 50835
rect 0 50663 624 50711
rect 330 50505 438 50615
rect 0 50409 624 50457
rect 330 50285 438 50361
rect 0 50189 624 50237
rect 0 50093 624 50141
rect 330 49969 438 50045
rect 0 49873 624 49921
rect 330 49715 438 49825
rect 0 49619 624 49667
rect 330 49495 438 49571
rect 0 49399 624 49447
rect 0 49303 624 49351
rect 330 49179 438 49255
rect 0 49083 624 49131
rect 330 48925 438 49035
rect 0 48829 624 48877
rect 330 48705 438 48781
rect 0 48609 624 48657
rect 0 48513 624 48561
rect 330 48389 438 48465
rect 0 48293 624 48341
rect 330 48135 438 48245
rect 0 48039 624 48087
rect 330 47915 438 47991
rect 0 47819 624 47867
rect 0 47723 624 47771
rect 330 47599 438 47675
rect 0 47503 624 47551
rect 330 47345 438 47455
rect 0 47249 624 47297
rect 330 47125 438 47201
rect 0 47029 624 47077
rect 0 46933 624 46981
rect 330 46809 438 46885
rect 0 46713 624 46761
rect 330 46555 438 46665
rect 0 46459 624 46507
rect 330 46335 438 46411
rect 0 46239 624 46287
rect 0 46143 624 46191
rect 330 46019 438 46095
rect 0 45923 624 45971
rect 330 45765 438 45875
rect 0 45669 624 45717
rect 330 45545 438 45621
rect 0 45449 624 45497
rect 0 45353 624 45401
rect 330 45229 438 45305
rect 0 45133 624 45181
rect 330 44975 438 45085
rect 0 44879 624 44927
rect 330 44755 438 44831
rect 0 44659 624 44707
rect 0 44563 624 44611
rect 330 44439 438 44515
rect 0 44343 624 44391
rect 330 44185 438 44295
rect 0 44089 624 44137
rect 330 43965 438 44041
rect 0 43869 624 43917
rect 0 43773 624 43821
rect 330 43649 438 43725
rect 0 43553 624 43601
rect 330 43395 438 43505
rect 0 43299 624 43347
rect 330 43175 438 43251
rect 0 43079 624 43127
rect 0 42983 624 43031
rect 330 42859 438 42935
rect 0 42763 624 42811
rect 330 42605 438 42715
rect 0 42509 624 42557
rect 330 42385 438 42461
rect 0 42289 624 42337
rect 0 42193 624 42241
rect 330 42069 438 42145
rect 0 41973 624 42021
rect 330 41815 438 41925
rect 0 41719 624 41767
rect 330 41595 438 41671
rect 0 41499 624 41547
rect 0 41403 624 41451
rect 330 41279 438 41355
rect 0 41183 624 41231
rect 330 41025 438 41135
rect 0 40929 624 40977
rect 330 40805 438 40881
rect 0 40709 624 40757
rect 0 40613 624 40661
rect 330 40489 438 40565
rect 0 40393 624 40441
rect 330 40235 438 40345
rect 0 40139 624 40187
rect 330 40015 438 40091
rect 0 39919 624 39967
rect 0 39823 624 39871
rect 330 39699 438 39775
rect 0 39603 624 39651
rect 330 39445 438 39555
rect 0 39349 624 39397
rect 330 39225 438 39301
rect 0 39129 624 39177
rect 0 39033 624 39081
rect 330 38909 438 38985
rect 0 38813 624 38861
rect 330 38655 438 38765
rect 0 38559 624 38607
rect 330 38435 438 38511
rect 0 38339 624 38387
rect 0 38243 624 38291
rect 330 38119 438 38195
rect 0 38023 624 38071
rect 330 37865 438 37975
rect 0 37769 624 37817
rect 330 37645 438 37721
rect 0 37549 624 37597
rect 0 37453 624 37501
rect 330 37329 438 37405
rect 0 37233 624 37281
rect 330 37075 438 37185
rect 0 36979 624 37027
rect 330 36855 438 36931
rect 0 36759 624 36807
rect 0 36663 624 36711
rect 330 36539 438 36615
rect 0 36443 624 36491
rect 330 36285 438 36395
rect 0 36189 624 36237
rect 330 36065 438 36141
rect 0 35969 624 36017
rect 0 35873 624 35921
rect 330 35749 438 35825
rect 0 35653 624 35701
rect 330 35495 438 35605
rect 0 35399 624 35447
rect 330 35275 438 35351
rect 0 35179 624 35227
rect 0 35083 624 35131
rect 330 34959 438 35035
rect 0 34863 624 34911
rect 330 34705 438 34815
rect 0 34609 624 34657
rect 330 34485 438 34561
rect 0 34389 624 34437
rect 0 34293 624 34341
rect 330 34169 438 34245
rect 0 34073 624 34121
rect 330 33915 438 34025
rect 0 33819 624 33867
rect 330 33695 438 33771
rect 0 33599 624 33647
rect 0 33503 624 33551
rect 330 33379 438 33455
rect 0 33283 624 33331
rect 330 33125 438 33235
rect 0 33029 624 33077
rect 330 32905 438 32981
rect 0 32809 624 32857
rect 0 32713 624 32761
rect 330 32589 438 32665
rect 0 32493 624 32541
rect 330 32335 438 32445
rect 0 32239 624 32287
rect 330 32115 438 32191
rect 0 32019 624 32067
rect 0 31923 624 31971
rect 330 31799 438 31875
rect 0 31703 624 31751
rect 330 31545 438 31655
rect 0 31449 624 31497
rect 330 31325 438 31401
rect 0 31229 624 31277
rect 0 31133 624 31181
rect 330 31009 438 31085
rect 0 30913 624 30961
rect 330 30755 438 30865
rect 0 30659 624 30707
rect 330 30535 438 30611
rect 0 30439 624 30487
rect 0 30343 624 30391
rect 330 30219 438 30295
rect 0 30123 624 30171
rect 330 29965 438 30075
rect 0 29869 624 29917
rect 330 29745 438 29821
rect 0 29649 624 29697
rect 0 29553 624 29601
rect 330 29429 438 29505
rect 0 29333 624 29381
rect 330 29175 438 29285
rect 0 29079 624 29127
rect 330 28955 438 29031
rect 0 28859 624 28907
rect 0 28763 624 28811
rect 330 28639 438 28715
rect 0 28543 624 28591
rect 330 28385 438 28495
rect 0 28289 624 28337
rect 330 28165 438 28241
rect 0 28069 624 28117
rect 0 27973 624 28021
rect 330 27849 438 27925
rect 0 27753 624 27801
rect 330 27595 438 27705
rect 0 27499 624 27547
rect 330 27375 438 27451
rect 0 27279 624 27327
rect 0 27183 624 27231
rect 330 27059 438 27135
rect 0 26963 624 27011
rect 330 26805 438 26915
rect 0 26709 624 26757
rect 330 26585 438 26661
rect 0 26489 624 26537
rect 0 26393 624 26441
rect 330 26269 438 26345
rect 0 26173 624 26221
rect 330 26015 438 26125
rect 0 25919 624 25967
rect 330 25795 438 25871
rect 0 25699 624 25747
rect 0 25603 624 25651
rect 330 25479 438 25555
rect 0 25383 624 25431
rect 330 25225 438 25335
rect 0 25129 624 25177
rect 330 25005 438 25081
rect 0 24909 624 24957
rect 0 24813 624 24861
rect 330 24689 438 24765
rect 0 24593 624 24641
rect 330 24435 438 24545
rect 0 24339 624 24387
rect 330 24215 438 24291
rect 0 24119 624 24167
rect 0 24023 624 24071
rect 330 23899 438 23975
rect 0 23803 624 23851
rect 330 23645 438 23755
rect 0 23549 624 23597
rect 330 23425 438 23501
rect 0 23329 624 23377
rect 0 23233 624 23281
rect 330 23109 438 23185
rect 0 23013 624 23061
rect 330 22855 438 22965
rect 0 22759 624 22807
rect 330 22635 438 22711
rect 0 22539 624 22587
rect 0 22443 624 22491
rect 330 22319 438 22395
rect 0 22223 624 22271
rect 330 22065 438 22175
rect 0 21969 624 22017
rect 330 21845 438 21921
rect 0 21749 624 21797
rect 0 21653 624 21701
rect 330 21529 438 21605
rect 0 21433 624 21481
rect 330 21275 438 21385
rect 0 21179 624 21227
rect 330 21055 438 21131
rect 0 20959 624 21007
rect 0 20863 624 20911
rect 330 20739 438 20815
rect 0 20643 624 20691
rect 330 20485 438 20595
rect 0 20389 624 20437
rect 330 20265 438 20341
rect 0 20169 624 20217
rect 0 20073 624 20121
rect 330 19949 438 20025
rect 0 19853 624 19901
rect 330 19695 438 19805
rect 0 19599 624 19647
rect 330 19475 438 19551
rect 0 19379 624 19427
rect 0 19283 624 19331
rect 330 19159 438 19235
rect 0 19063 624 19111
rect 330 18905 438 19015
rect 0 18809 624 18857
rect 330 18685 438 18761
rect 0 18589 624 18637
rect 0 18493 624 18541
rect 330 18369 438 18445
rect 0 18273 624 18321
rect 330 18115 438 18225
rect 0 18019 624 18067
rect 330 17895 438 17971
rect 0 17799 624 17847
rect 0 17703 624 17751
rect 330 17579 438 17655
rect 0 17483 624 17531
rect 330 17325 438 17435
rect 0 17229 624 17277
rect 330 17105 438 17181
rect 0 17009 624 17057
rect 0 16913 624 16961
rect 330 16789 438 16865
rect 0 16693 624 16741
rect 330 16535 438 16645
rect 0 16439 624 16487
rect 330 16315 438 16391
rect 0 16219 624 16267
rect 0 16123 624 16171
rect 330 15999 438 16075
rect 0 15903 624 15951
rect 330 15745 438 15855
rect 0 15649 624 15697
rect 330 15525 438 15601
rect 0 15429 624 15477
rect 0 15333 624 15381
rect 330 15209 438 15285
rect 0 15113 624 15161
rect 330 14955 438 15065
rect 0 14859 624 14907
rect 330 14735 438 14811
rect 0 14639 624 14687
rect 0 14543 624 14591
rect 330 14419 438 14495
rect 0 14323 624 14371
rect 330 14165 438 14275
rect 0 14069 624 14117
rect 330 13945 438 14021
rect 0 13849 624 13897
rect 0 13753 624 13801
rect 330 13629 438 13705
rect 0 13533 624 13581
rect 330 13375 438 13485
rect 0 13279 624 13327
rect 330 13155 438 13231
rect 0 13059 624 13107
rect 0 12963 624 13011
rect 330 12839 438 12915
rect 0 12743 624 12791
rect 330 12585 438 12695
rect 0 12489 624 12537
rect 330 12365 438 12441
rect 0 12269 624 12317
rect 0 12173 624 12221
rect 330 12049 438 12125
rect 0 11953 624 12001
rect 330 11795 438 11905
rect 0 11699 624 11747
rect 330 11575 438 11651
rect 0 11479 624 11527
rect 0 11383 624 11431
rect 330 11259 438 11335
rect 0 11163 624 11211
rect 330 11005 438 11115
rect 0 10909 624 10957
rect 330 10785 438 10861
rect 0 10689 624 10737
rect 0 10593 624 10641
rect 330 10469 438 10545
rect 0 10373 624 10421
rect 330 10215 438 10325
rect 0 10119 624 10167
rect 330 9995 438 10071
rect 0 9899 624 9947
rect 0 9803 624 9851
rect 330 9679 438 9755
rect 0 9583 624 9631
rect 330 9425 438 9535
rect 0 9329 624 9377
rect 330 9205 438 9281
rect 0 9109 624 9157
rect 0 9013 624 9061
rect 330 8889 438 8965
rect 0 8793 624 8841
rect 330 8635 438 8745
rect 0 8539 624 8587
rect 330 8415 438 8491
rect 0 8319 624 8367
rect 0 8223 624 8271
rect 330 8099 438 8175
rect 0 8003 624 8051
rect 330 7845 438 7955
rect 0 7749 624 7797
rect 330 7625 438 7701
rect 0 7529 624 7577
rect 0 7433 624 7481
rect 330 7309 438 7385
rect 0 7213 624 7261
rect 330 7055 438 7165
rect 0 6959 624 7007
rect 330 6835 438 6911
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 330 6519 438 6595
rect 0 6423 624 6471
rect 330 6265 438 6375
rect 0 6169 624 6217
rect 330 6045 438 6121
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 330 5729 438 5805
rect 0 5633 624 5681
rect 330 5475 438 5585
rect 0 5379 624 5427
rect 330 5255 438 5331
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 330 4939 438 5015
rect 0 4843 624 4891
rect 330 4685 438 4795
rect 0 4589 624 4637
rect 330 4465 438 4541
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 330 4149 438 4225
rect 0 4053 624 4101
rect 330 3895 438 4005
rect 0 3799 624 3847
rect 330 3675 438 3751
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 330 3359 438 3435
rect 0 3263 624 3311
rect 330 3105 438 3215
rect 0 3009 624 3057
rect 330 2885 438 2961
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 330 2569 438 2645
rect 0 2473 624 2521
rect 330 2315 438 2425
rect 0 2219 624 2267
rect 330 2095 438 2171
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 330 1779 438 1855
rect 0 1683 624 1731
rect 330 1525 438 1635
rect 0 1429 624 1477
rect 330 1305 438 1381
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 330 989 438 1065
rect 0 893 624 941
rect 330 735 438 845
rect 0 639 624 687
rect 330 515 438 591
rect 0 419 624 467
rect 284 257 340 266
rect 284 192 340 201
<< via2 >>
rect 284 51883 340 51939
rect 284 201 340 257
<< metal3 >>
rect 263 51939 361 51960
rect 263 51883 284 51939
rect 340 51883 361 51939
rect 263 51862 361 51883
rect 263 257 361 278
rect 263 201 284 257
rect 340 201 361 257
rect 263 180 361 201
use sky130_fd_bd_sram__openram_dp_cell_cap_col_3  sky130_fd_bd_sram__openram_dp_cell_cap_col_0
timestamp 1676037725
transform -1 0 624 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col_3  sky130_fd_bd_sram__openram_dp_cell_cap_col_1
timestamp 1676037725
transform -1 0 624 0 -1 52140
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_dummy_3  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1676037725
transform -1 0 624 0 1 51350
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_0
timestamp 1676037725
transform -1 0 624 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_1
timestamp 1676037725
transform -1 0 624 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_2
timestamp 1676037725
transform -1 0 624 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_3
timestamp 1676037725
transform -1 0 624 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_4
timestamp 1676037725
transform -1 0 624 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_5
timestamp 1676037725
transform -1 0 624 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_6
timestamp 1676037725
transform -1 0 624 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_7
timestamp 1676037725
transform -1 0 624 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_8
timestamp 1676037725
transform -1 0 624 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_9
timestamp 1676037725
transform -1 0 624 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_10
timestamp 1676037725
transform -1 0 624 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_11
timestamp 1676037725
transform -1 0 624 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_12
timestamp 1676037725
transform -1 0 624 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_13
timestamp 1676037725
transform -1 0 624 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_14
timestamp 1676037725
transform -1 0 624 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_15
timestamp 1676037725
transform -1 0 624 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_16
timestamp 1676037725
transform -1 0 624 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_17
timestamp 1676037725
transform -1 0 624 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_18
timestamp 1676037725
transform -1 0 624 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_19
timestamp 1676037725
transform -1 0 624 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_20
timestamp 1676037725
transform -1 0 624 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_21
timestamp 1676037725
transform -1 0 624 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_22
timestamp 1676037725
transform -1 0 624 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_23
timestamp 1676037725
transform -1 0 624 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_24
timestamp 1676037725
transform -1 0 624 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_25
timestamp 1676037725
transform -1 0 624 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_26
timestamp 1676037725
transform -1 0 624 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_27
timestamp 1676037725
transform -1 0 624 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_28
timestamp 1676037725
transform -1 0 624 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_29
timestamp 1676037725
transform -1 0 624 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_30
timestamp 1676037725
transform -1 0 624 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_31
timestamp 1676037725
transform -1 0 624 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_32
timestamp 1676037725
transform -1 0 624 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_33
timestamp 1676037725
transform -1 0 624 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_34
timestamp 1676037725
transform -1 0 624 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_35
timestamp 1676037725
transform -1 0 624 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_36
timestamp 1676037725
transform -1 0 624 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_37
timestamp 1676037725
transform -1 0 624 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_38
timestamp 1676037725
transform -1 0 624 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_39
timestamp 1676037725
transform -1 0 624 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_40
timestamp 1676037725
transform -1 0 624 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_41
timestamp 1676037725
transform -1 0 624 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_42
timestamp 1676037725
transform -1 0 624 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_43
timestamp 1676037725
transform -1 0 624 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_44
timestamp 1676037725
transform -1 0 624 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_45
timestamp 1676037725
transform -1 0 624 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_46
timestamp 1676037725
transform -1 0 624 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_47
timestamp 1676037725
transform -1 0 624 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_48
timestamp 1676037725
transform -1 0 624 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_49
timestamp 1676037725
transform -1 0 624 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_50
timestamp 1676037725
transform -1 0 624 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_51
timestamp 1676037725
transform -1 0 624 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_52
timestamp 1676037725
transform -1 0 624 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_53
timestamp 1676037725
transform -1 0 624 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_54
timestamp 1676037725
transform -1 0 624 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_55
timestamp 1676037725
transform -1 0 624 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_56
timestamp 1676037725
transform -1 0 624 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_57
timestamp 1676037725
transform -1 0 624 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_58
timestamp 1676037725
transform -1 0 624 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_59
timestamp 1676037725
transform -1 0 624 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_60
timestamp 1676037725
transform -1 0 624 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_61
timestamp 1676037725
transform -1 0 624 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_62
timestamp 1676037725
transform -1 0 624 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_63
timestamp 1676037725
transform -1 0 624 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_64
timestamp 1676037725
transform -1 0 624 0 -1 51350
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_65
timestamp 1676037725
transform -1 0 624 0 1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_66
timestamp 1676037725
transform -1 0 624 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_67
timestamp 1676037725
transform -1 0 624 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_68
timestamp 1676037725
transform -1 0 624 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_69
timestamp 1676037725
transform -1 0 624 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_70
timestamp 1676037725
transform -1 0 624 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_71
timestamp 1676037725
transform -1 0 624 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_72
timestamp 1676037725
transform -1 0 624 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_73
timestamp 1676037725
transform -1 0 624 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_74
timestamp 1676037725
transform -1 0 624 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_75
timestamp 1676037725
transform -1 0 624 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_76
timestamp 1676037725
transform -1 0 624 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_77
timestamp 1676037725
transform -1 0 624 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_78
timestamp 1676037725
transform -1 0 624 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_79
timestamp 1676037725
transform -1 0 624 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_80
timestamp 1676037725
transform -1 0 624 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_81
timestamp 1676037725
transform -1 0 624 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_82
timestamp 1676037725
transform -1 0 624 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_83
timestamp 1676037725
transform -1 0 624 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_84
timestamp 1676037725
transform -1 0 624 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_85
timestamp 1676037725
transform -1 0 624 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_86
timestamp 1676037725
transform -1 0 624 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_87
timestamp 1676037725
transform -1 0 624 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_88
timestamp 1676037725
transform -1 0 624 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_89
timestamp 1676037725
transform -1 0 624 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_90
timestamp 1676037725
transform -1 0 624 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_91
timestamp 1676037725
transform -1 0 624 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_92
timestamp 1676037725
transform -1 0 624 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_93
timestamp 1676037725
transform -1 0 624 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_94
timestamp 1676037725
transform -1 0 624 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_95
timestamp 1676037725
transform -1 0 624 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_96
timestamp 1676037725
transform -1 0 624 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_97
timestamp 1676037725
transform -1 0 624 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_98
timestamp 1676037725
transform -1 0 624 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_99
timestamp 1676037725
transform -1 0 624 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_100
timestamp 1676037725
transform -1 0 624 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_101
timestamp 1676037725
transform -1 0 624 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_102
timestamp 1676037725
transform -1 0 624 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_103
timestamp 1676037725
transform -1 0 624 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_104
timestamp 1676037725
transform -1 0 624 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_105
timestamp 1676037725
transform -1 0 624 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_106
timestamp 1676037725
transform -1 0 624 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_107
timestamp 1676037725
transform -1 0 624 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_108
timestamp 1676037725
transform -1 0 624 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_109
timestamp 1676037725
transform -1 0 624 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_110
timestamp 1676037725
transform -1 0 624 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_111
timestamp 1676037725
transform -1 0 624 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_112
timestamp 1676037725
transform -1 0 624 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_113
timestamp 1676037725
transform -1 0 624 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_114
timestamp 1676037725
transform -1 0 624 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_115
timestamp 1676037725
transform -1 0 624 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_116
timestamp 1676037725
transform -1 0 624 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_117
timestamp 1676037725
transform -1 0 624 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_118
timestamp 1676037725
transform -1 0 624 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_119
timestamp 1676037725
transform -1 0 624 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_120
timestamp 1676037725
transform -1 0 624 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_121
timestamp 1676037725
transform -1 0 624 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_122
timestamp 1676037725
transform -1 0 624 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_123
timestamp 1676037725
transform -1 0 624 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_124
timestamp 1676037725
transform -1 0 624 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_125
timestamp 1676037725
transform -1 0 624 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_126
timestamp 1676037725
transform -1 0 624 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_127
timestamp 1676037725
transform -1 0 624 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_3  sky130_fd_bd_sram__openram_dp_cell_replica_128
timestamp 1676037725
transform -1 0 624 0 -1 26070
box -42 -105 650 421
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_0
timestamp 1676037725
transform 1 0 279 0 1 192
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_1
timestamp 1676037725
transform 1 0 279 0 1 51874
box 0 0 1 1
<< labels >>
rlabel metal3 s 263 51862 361 51960 4 vdd
rlabel metal3 s 263 180 361 278 4 vdd
rlabel metal2 s 330 50759 438 50835 4 gnd
rlabel metal2 s 330 48135 438 48245 4 gnd
rlabel metal2 s 330 36539 438 36615 4 gnd
rlabel metal2 s 330 28385 438 28495 4 gnd
rlabel metal2 s 330 51295 438 51405 4 gnd
rlabel metal2 s 330 41815 438 41925 4 gnd
rlabel metal2 s 330 29175 438 29285 4 gnd
rlabel metal2 s 330 30219 438 30295 4 gnd
rlabel metal2 s 330 36065 438 36141 4 gnd
rlabel metal2 s 330 50285 438 50361 4 gnd
rlabel metal2 s 330 34705 438 34815 4 gnd
rlabel metal2 s 330 43649 438 43725 4 gnd
rlabel metal2 s 330 28955 438 29031 4 gnd
rlabel metal2 s 330 45229 438 45305 4 gnd
rlabel metal2 s 330 32115 438 32191 4 gnd
rlabel metal2 s 330 34485 438 34561 4 gnd
rlabel metal2 s 330 46019 438 46095 4 gnd
rlabel metal2 s 330 33695 438 33771 4 gnd
rlabel metal2 s 330 26269 438 26345 4 gnd
rlabel metal2 s 330 32589 438 32665 4 gnd
rlabel metal2 s 330 47345 438 47455 4 gnd
rlabel metal2 s 330 37865 438 37975 4 gnd
rlabel metal2 s 330 31325 438 31401 4 gnd
rlabel metal2 s 330 35749 438 35825 4 gnd
rlabel metal2 s 330 33125 438 33235 4 gnd
rlabel metal2 s 330 34959 438 35035 4 gnd
rlabel metal2 s 330 42385 438 42461 4 gnd
rlabel metal2 s 330 41279 438 41355 4 gnd
rlabel metal2 s 330 45545 438 45621 4 gnd
rlabel metal2 s 330 47599 438 47675 4 gnd
rlabel metal2 s 330 41025 438 41135 4 gnd
rlabel metal2 s 330 40489 438 40565 4 gnd
rlabel metal2 s 330 43965 438 44041 4 gnd
rlabel metal2 s 330 28165 438 28241 4 gnd
rlabel metal2 s 330 43395 438 43505 4 gnd
rlabel metal2 s 330 31545 438 31655 4 gnd
rlabel metal2 s 330 38119 438 38195 4 gnd
rlabel metal2 s 330 39445 438 39555 4 gnd
rlabel metal2 s 330 31009 438 31085 4 gnd
rlabel metal2 s 330 34169 438 34245 4 gnd
rlabel metal2 s 330 50505 438 50615 4 gnd
rlabel metal2 s 330 42859 438 42935 4 gnd
rlabel metal2 s 330 27595 438 27705 4 gnd
rlabel metal2 s 330 27849 438 27925 4 gnd
rlabel metal2 s 330 35275 438 35351 4 gnd
rlabel metal2 s 330 41595 438 41671 4 gnd
rlabel metal2 s 330 51075 438 51151 4 gnd
rlabel metal2 s 330 39225 438 39301 4 gnd
rlabel metal2 s 330 46555 438 46665 4 gnd
rlabel metal2 s 330 37329 438 37405 4 gnd
rlabel metal2 s 330 40235 438 40345 4 gnd
rlabel metal2 s 330 49969 438 50045 4 gnd
rlabel metal2 s 330 33915 438 34025 4 gnd
rlabel metal2 s 330 40015 438 40091 4 gnd
rlabel metal2 s 330 44755 438 44831 4 gnd
rlabel metal2 s 330 38655 438 38765 4 gnd
rlabel metal2 s 330 48389 438 48465 4 gnd
rlabel metal2 s 330 33379 438 33455 4 gnd
rlabel metal2 s 330 44439 438 44515 4 gnd
rlabel metal2 s 330 27059 438 27135 4 gnd
rlabel metal2 s 330 32335 438 32445 4 gnd
rlabel metal2 s 330 42069 438 42145 4 gnd
rlabel metal2 s 330 45765 438 45875 4 gnd
rlabel metal2 s 330 36855 438 36931 4 gnd
rlabel metal2 s 330 49715 438 49825 4 gnd
rlabel metal2 s 330 51549 438 51625 4 gnd
rlabel metal2 s 330 37075 438 37185 4 gnd
rlabel metal2 s 330 37645 438 37721 4 gnd
rlabel metal2 s 330 26585 438 26661 4 gnd
rlabel metal2 s 330 40805 438 40881 4 gnd
rlabel metal2 s 330 39699 438 39775 4 gnd
rlabel metal2 s 330 35495 438 35605 4 gnd
rlabel metal2 s 330 30535 438 30611 4 gnd
rlabel metal2 s 330 47125 438 47201 4 gnd
rlabel metal2 s 330 26805 438 26915 4 gnd
rlabel metal2 s 330 31799 438 31875 4 gnd
rlabel metal2 s 330 27375 438 27451 4 gnd
rlabel metal2 s 330 38909 438 38985 4 gnd
rlabel metal2 s 330 44185 438 44295 4 gnd
rlabel metal2 s 330 42605 438 42715 4 gnd
rlabel metal2 s 330 38435 438 38511 4 gnd
rlabel metal2 s 330 46809 438 46885 4 gnd
rlabel metal2 s 330 48705 438 48781 4 gnd
rlabel metal2 s 330 30755 438 30865 4 gnd
rlabel metal2 s 330 47915 438 47991 4 gnd
rlabel metal2 s 330 43175 438 43251 4 gnd
rlabel metal2 s 330 44975 438 45085 4 gnd
rlabel metal2 s 330 28639 438 28715 4 gnd
rlabel metal2 s 330 36285 438 36395 4 gnd
rlabel metal2 s 330 29965 438 30075 4 gnd
rlabel metal2 s 330 29429 438 29505 4 gnd
rlabel metal2 s 330 49179 438 49255 4 gnd
rlabel metal2 s 330 29745 438 29821 4 gnd
rlabel metal2 s 330 32905 438 32981 4 gnd
rlabel metal2 s 330 48925 438 49035 4 gnd
rlabel metal2 s 330 46335 438 46411 4 gnd
rlabel metal2 s 330 49495 438 49571 4 gnd
rlabel metal2 s 0 39349 624 39397 4 wl_1_98
rlabel metal2 s 0 39603 624 39651 4 wl_1_99
rlabel metal2 s 0 40139 624 40187 4 wl_1_100
rlabel metal2 s 0 40393 624 40441 4 wl_1_101
rlabel metal2 s 0 40929 624 40977 4 wl_1_102
rlabel metal2 s 0 41183 624 41231 4 wl_1_103
rlabel metal2 s 0 41719 624 41767 4 wl_1_104
rlabel metal2 s 0 41973 624 42021 4 wl_1_105
rlabel metal2 s 0 42509 624 42557 4 wl_1_106
rlabel metal2 s 0 42763 624 42811 4 wl_1_107
rlabel metal2 s 0 43299 624 43347 4 wl_1_108
rlabel metal2 s 0 43553 624 43601 4 wl_1_109
rlabel metal2 s 0 44089 624 44137 4 wl_1_110
rlabel metal2 s 0 44343 624 44391 4 wl_1_111
rlabel metal2 s 0 44879 624 44927 4 wl_1_112
rlabel metal2 s 0 45133 624 45181 4 wl_1_113
rlabel metal2 s 0 45669 624 45717 4 wl_1_114
rlabel metal2 s 0 45923 624 45971 4 wl_1_115
rlabel metal2 s 0 46459 624 46507 4 wl_1_116
rlabel metal2 s 0 46713 624 46761 4 wl_1_117
rlabel metal2 s 0 47249 624 47297 4 wl_1_118
rlabel metal2 s 0 47503 624 47551 4 wl_1_119
rlabel metal2 s 0 48039 624 48087 4 wl_1_120
rlabel metal2 s 0 48293 624 48341 4 wl_1_121
rlabel metal2 s 0 48829 624 48877 4 wl_1_122
rlabel metal2 s 0 49083 624 49131 4 wl_1_123
rlabel metal2 s 0 49619 624 49667 4 wl_1_124
rlabel metal2 s 0 49873 624 49921 4 wl_1_125
rlabel metal2 s 0 50409 624 50457 4 wl_1_126
rlabel metal2 s 0 50663 624 50711 4 wl_1_127
rlabel metal2 s 0 51199 624 51247 4 wl_1_128
rlabel metal2 s 0 51453 624 51501 4 wl_1_129
rlabel metal2 s 0 39033 624 39081 4 wl_0_97
rlabel metal2 s 0 39129 624 39177 4 wl_0_98
rlabel metal2 s 0 39823 624 39871 4 wl_0_99
rlabel metal2 s 0 39919 624 39967 4 wl_0_100
rlabel metal2 s 0 40613 624 40661 4 wl_0_101
rlabel metal2 s 0 40709 624 40757 4 wl_0_102
rlabel metal2 s 0 41403 624 41451 4 wl_0_103
rlabel metal2 s 0 41499 624 41547 4 wl_0_104
rlabel metal2 s 0 42193 624 42241 4 wl_0_105
rlabel metal2 s 0 42289 624 42337 4 wl_0_106
rlabel metal2 s 0 42983 624 43031 4 wl_0_107
rlabel metal2 s 0 43079 624 43127 4 wl_0_108
rlabel metal2 s 0 43773 624 43821 4 wl_0_109
rlabel metal2 s 0 43869 624 43917 4 wl_0_110
rlabel metal2 s 0 44563 624 44611 4 wl_0_111
rlabel metal2 s 0 44659 624 44707 4 wl_0_112
rlabel metal2 s 0 45353 624 45401 4 wl_0_113
rlabel metal2 s 0 45449 624 45497 4 wl_0_114
rlabel metal2 s 0 46143 624 46191 4 wl_0_115
rlabel metal2 s 0 46239 624 46287 4 wl_0_116
rlabel metal2 s 0 46933 624 46981 4 wl_0_117
rlabel metal2 s 0 47029 624 47077 4 wl_0_118
rlabel metal2 s 0 47723 624 47771 4 wl_0_119
rlabel metal2 s 0 47819 624 47867 4 wl_0_120
rlabel metal2 s 0 48513 624 48561 4 wl_0_121
rlabel metal2 s 0 48609 624 48657 4 wl_0_122
rlabel metal2 s 0 49303 624 49351 4 wl_0_123
rlabel metal2 s 0 49399 624 49447 4 wl_0_124
rlabel metal2 s 0 50093 624 50141 4 wl_0_125
rlabel metal2 s 0 50189 624 50237 4 wl_0_126
rlabel metal2 s 0 50883 624 50931 4 wl_0_127
rlabel metal2 s 0 50979 624 51027 4 wl_0_128
rlabel metal2 s 0 51673 624 51721 4 wl_0_129
rlabel metal2 s 0 38813 624 38861 4 wl_1_97
rlabel metal2 s 0 26393 624 26441 4 wl_0_65
rlabel metal2 s 0 26489 624 26537 4 wl_0_66
rlabel metal2 s 0 27183 624 27231 4 wl_0_67
rlabel metal2 s 0 27279 624 27327 4 wl_0_68
rlabel metal2 s 0 27973 624 28021 4 wl_0_69
rlabel metal2 s 0 28069 624 28117 4 wl_0_70
rlabel metal2 s 0 28763 624 28811 4 wl_0_71
rlabel metal2 s 0 28859 624 28907 4 wl_0_72
rlabel metal2 s 0 29553 624 29601 4 wl_0_73
rlabel metal2 s 0 29649 624 29697 4 wl_0_74
rlabel metal2 s 0 30343 624 30391 4 wl_0_75
rlabel metal2 s 0 30439 624 30487 4 wl_0_76
rlabel metal2 s 0 31133 624 31181 4 wl_0_77
rlabel metal2 s 0 31229 624 31277 4 wl_0_78
rlabel metal2 s 0 31923 624 31971 4 wl_0_79
rlabel metal2 s 0 32019 624 32067 4 wl_0_80
rlabel metal2 s 0 32713 624 32761 4 wl_0_81
rlabel metal2 s 0 32809 624 32857 4 wl_0_82
rlabel metal2 s 0 33503 624 33551 4 wl_0_83
rlabel metal2 s 0 33599 624 33647 4 wl_0_84
rlabel metal2 s 0 34293 624 34341 4 wl_0_85
rlabel metal2 s 0 34389 624 34437 4 wl_0_86
rlabel metal2 s 0 35083 624 35131 4 wl_0_87
rlabel metal2 s 0 35179 624 35227 4 wl_0_88
rlabel metal2 s 0 35873 624 35921 4 wl_0_89
rlabel metal2 s 0 35969 624 36017 4 wl_0_90
rlabel metal2 s 0 36663 624 36711 4 wl_0_91
rlabel metal2 s 0 36759 624 36807 4 wl_0_92
rlabel metal2 s 0 37453 624 37501 4 wl_0_93
rlabel metal2 s 0 37549 624 37597 4 wl_0_94
rlabel metal2 s 0 38243 624 38291 4 wl_0_95
rlabel metal2 s 0 38339 624 38387 4 wl_0_96
rlabel metal2 s 0 26173 624 26221 4 wl_1_65
rlabel metal2 s 0 26709 624 26757 4 wl_1_66
rlabel metal2 s 0 26963 624 27011 4 wl_1_67
rlabel metal2 s 0 27499 624 27547 4 wl_1_68
rlabel metal2 s 0 27753 624 27801 4 wl_1_69
rlabel metal2 s 0 28289 624 28337 4 wl_1_70
rlabel metal2 s 0 28543 624 28591 4 wl_1_71
rlabel metal2 s 0 29079 624 29127 4 wl_1_72
rlabel metal2 s 0 29333 624 29381 4 wl_1_73
rlabel metal2 s 0 29869 624 29917 4 wl_1_74
rlabel metal2 s 0 30123 624 30171 4 wl_1_75
rlabel metal2 s 0 30659 624 30707 4 wl_1_76
rlabel metal2 s 0 30913 624 30961 4 wl_1_77
rlabel metal2 s 0 31449 624 31497 4 wl_1_78
rlabel metal2 s 0 31703 624 31751 4 wl_1_79
rlabel metal2 s 0 32239 624 32287 4 wl_1_80
rlabel metal2 s 0 32493 624 32541 4 wl_1_81
rlabel metal2 s 0 33029 624 33077 4 wl_1_82
rlabel metal2 s 0 33283 624 33331 4 wl_1_83
rlabel metal2 s 0 33819 624 33867 4 wl_1_84
rlabel metal2 s 0 34073 624 34121 4 wl_1_85
rlabel metal2 s 0 34609 624 34657 4 wl_1_86
rlabel metal2 s 0 34863 624 34911 4 wl_1_87
rlabel metal2 s 0 35399 624 35447 4 wl_1_88
rlabel metal2 s 0 35653 624 35701 4 wl_1_89
rlabel metal2 s 0 36189 624 36237 4 wl_1_90
rlabel metal2 s 0 36443 624 36491 4 wl_1_91
rlabel metal2 s 0 36979 624 37027 4 wl_1_92
rlabel metal2 s 0 37233 624 37281 4 wl_1_93
rlabel metal2 s 0 37769 624 37817 4 wl_1_94
rlabel metal2 s 0 38023 624 38071 4 wl_1_95
rlabel metal2 s 0 38559 624 38607 4 wl_1_96
rlabel metal2 s 0 13753 624 13801 4 wl_0_33
rlabel metal2 s 0 13849 624 13897 4 wl_0_34
rlabel metal2 s 0 14543 624 14591 4 wl_0_35
rlabel metal2 s 0 14639 624 14687 4 wl_0_36
rlabel metal2 s 0 15333 624 15381 4 wl_0_37
rlabel metal2 s 0 15429 624 15477 4 wl_0_38
rlabel metal2 s 0 16123 624 16171 4 wl_0_39
rlabel metal2 s 0 16219 624 16267 4 wl_0_40
rlabel metal2 s 0 16913 624 16961 4 wl_0_41
rlabel metal2 s 0 17009 624 17057 4 wl_0_42
rlabel metal2 s 0 17703 624 17751 4 wl_0_43
rlabel metal2 s 0 17799 624 17847 4 wl_0_44
rlabel metal2 s 0 18493 624 18541 4 wl_0_45
rlabel metal2 s 0 18589 624 18637 4 wl_0_46
rlabel metal2 s 0 19283 624 19331 4 wl_0_47
rlabel metal2 s 0 19379 624 19427 4 wl_0_48
rlabel metal2 s 0 20073 624 20121 4 wl_0_49
rlabel metal2 s 0 20169 624 20217 4 wl_0_50
rlabel metal2 s 0 20863 624 20911 4 wl_0_51
rlabel metal2 s 0 20959 624 21007 4 wl_0_52
rlabel metal2 s 0 21653 624 21701 4 wl_0_53
rlabel metal2 s 0 21749 624 21797 4 wl_0_54
rlabel metal2 s 0 22443 624 22491 4 wl_0_55
rlabel metal2 s 0 22539 624 22587 4 wl_0_56
rlabel metal2 s 0 23233 624 23281 4 wl_0_57
rlabel metal2 s 0 23329 624 23377 4 wl_0_58
rlabel metal2 s 0 24023 624 24071 4 wl_0_59
rlabel metal2 s 0 24119 624 24167 4 wl_0_60
rlabel metal2 s 0 24813 624 24861 4 wl_0_61
rlabel metal2 s 0 24909 624 24957 4 wl_0_62
rlabel metal2 s 0 25603 624 25651 4 wl_0_63
rlabel metal2 s 0 25699 624 25747 4 wl_0_64
rlabel metal2 s 0 13279 624 13327 4 wl_1_32
rlabel metal2 s 0 13533 624 13581 4 wl_1_33
rlabel metal2 s 0 14069 624 14117 4 wl_1_34
rlabel metal2 s 0 14323 624 14371 4 wl_1_35
rlabel metal2 s 0 14859 624 14907 4 wl_1_36
rlabel metal2 s 0 15113 624 15161 4 wl_1_37
rlabel metal2 s 0 15649 624 15697 4 wl_1_38
rlabel metal2 s 0 15903 624 15951 4 wl_1_39
rlabel metal2 s 0 16439 624 16487 4 wl_1_40
rlabel metal2 s 0 16693 624 16741 4 wl_1_41
rlabel metal2 s 0 17229 624 17277 4 wl_1_42
rlabel metal2 s 0 17483 624 17531 4 wl_1_43
rlabel metal2 s 0 18019 624 18067 4 wl_1_44
rlabel metal2 s 0 18273 624 18321 4 wl_1_45
rlabel metal2 s 0 18809 624 18857 4 wl_1_46
rlabel metal2 s 0 19063 624 19111 4 wl_1_47
rlabel metal2 s 0 19599 624 19647 4 wl_1_48
rlabel metal2 s 0 19853 624 19901 4 wl_1_49
rlabel metal2 s 0 20389 624 20437 4 wl_1_50
rlabel metal2 s 0 20643 624 20691 4 wl_1_51
rlabel metal2 s 0 21179 624 21227 4 wl_1_52
rlabel metal2 s 0 21433 624 21481 4 wl_1_53
rlabel metal2 s 0 21969 624 22017 4 wl_1_54
rlabel metal2 s 0 22223 624 22271 4 wl_1_55
rlabel metal2 s 0 22759 624 22807 4 wl_1_56
rlabel metal2 s 0 23013 624 23061 4 wl_1_57
rlabel metal2 s 0 23549 624 23597 4 wl_1_58
rlabel metal2 s 0 23803 624 23851 4 wl_1_59
rlabel metal2 s 0 24339 624 24387 4 wl_1_60
rlabel metal2 s 0 24593 624 24641 4 wl_1_61
rlabel metal2 s 0 25129 624 25177 4 wl_1_62
rlabel metal2 s 0 25383 624 25431 4 wl_1_63
rlabel metal2 s 0 25919 624 25967 4 wl_1_64
rlabel metal2 s 0 13059 624 13107 4 wl_0_32
rlabel metal2 s 0 639 624 687 4 wl_1_0
rlabel metal2 s 0 893 624 941 4 wl_1_1
rlabel metal2 s 0 1429 624 1477 4 wl_1_2
rlabel metal2 s 0 1683 624 1731 4 wl_1_3
rlabel metal2 s 0 2219 624 2267 4 wl_1_4
rlabel metal2 s 0 2473 624 2521 4 wl_1_5
rlabel metal2 s 0 3009 624 3057 4 wl_1_6
rlabel metal2 s 0 3263 624 3311 4 wl_1_7
rlabel metal2 s 0 3799 624 3847 4 wl_1_8
rlabel metal2 s 0 4053 624 4101 4 wl_1_9
rlabel metal2 s 0 4589 624 4637 4 wl_1_10
rlabel metal2 s 0 4843 624 4891 4 wl_1_11
rlabel metal2 s 0 5379 624 5427 4 wl_1_12
rlabel metal2 s 0 5633 624 5681 4 wl_1_13
rlabel metal2 s 0 6169 624 6217 4 wl_1_14
rlabel metal2 s 0 6423 624 6471 4 wl_1_15
rlabel metal2 s 0 6959 624 7007 4 wl_1_16
rlabel metal2 s 0 7213 624 7261 4 wl_1_17
rlabel metal2 s 0 7749 624 7797 4 wl_1_18
rlabel metal2 s 0 8003 624 8051 4 wl_1_19
rlabel metal2 s 0 8539 624 8587 4 wl_1_20
rlabel metal2 s 0 8793 624 8841 4 wl_1_21
rlabel metal2 s 0 9329 624 9377 4 wl_1_22
rlabel metal2 s 0 9583 624 9631 4 wl_1_23
rlabel metal2 s 0 10119 624 10167 4 wl_1_24
rlabel metal2 s 0 10373 624 10421 4 wl_1_25
rlabel metal2 s 0 10909 624 10957 4 wl_1_26
rlabel metal2 s 0 11163 624 11211 4 wl_1_27
rlabel metal2 s 0 11699 624 11747 4 wl_1_28
rlabel metal2 s 0 11953 624 12001 4 wl_1_29
rlabel metal2 s 0 12489 624 12537 4 wl_1_30
rlabel metal2 s 0 12743 624 12791 4 wl_1_31
rlabel metal2 s 0 419 624 467 4 wl_0_0
rlabel metal2 s 0 1113 624 1161 4 wl_0_1
rlabel metal2 s 0 1209 624 1257 4 wl_0_2
rlabel metal2 s 0 1903 624 1951 4 wl_0_3
rlabel metal2 s 0 1999 624 2047 4 wl_0_4
rlabel metal2 s 0 2693 624 2741 4 wl_0_5
rlabel metal2 s 0 2789 624 2837 4 wl_0_6
rlabel metal2 s 0 3483 624 3531 4 wl_0_7
rlabel metal2 s 0 3579 624 3627 4 wl_0_8
rlabel metal2 s 0 4273 624 4321 4 wl_0_9
rlabel metal2 s 0 4369 624 4417 4 wl_0_10
rlabel metal2 s 0 5063 624 5111 4 wl_0_11
rlabel metal2 s 0 5159 624 5207 4 wl_0_12
rlabel metal2 s 0 5853 624 5901 4 wl_0_13
rlabel metal2 s 0 5949 624 5997 4 wl_0_14
rlabel metal2 s 0 6643 624 6691 4 wl_0_15
rlabel metal2 s 0 6739 624 6787 4 wl_0_16
rlabel metal2 s 0 7433 624 7481 4 wl_0_17
rlabel metal2 s 0 7529 624 7577 4 wl_0_18
rlabel metal2 s 0 8223 624 8271 4 wl_0_19
rlabel metal2 s 0 8319 624 8367 4 wl_0_20
rlabel metal2 s 0 9013 624 9061 4 wl_0_21
rlabel metal2 s 0 9109 624 9157 4 wl_0_22
rlabel metal2 s 0 9803 624 9851 4 wl_0_23
rlabel metal2 s 0 9899 624 9947 4 wl_0_24
rlabel metal2 s 0 10593 624 10641 4 wl_0_25
rlabel metal2 s 0 10689 624 10737 4 wl_0_26
rlabel metal2 s 0 11383 624 11431 4 wl_0_27
rlabel metal2 s 0 11479 624 11527 4 wl_0_28
rlabel metal2 s 0 12173 624 12221 4 wl_0_29
rlabel metal2 s 0 12269 624 12317 4 wl_0_30
rlabel metal2 s 0 12963 624 13011 4 wl_0_31
rlabel metal2 s 330 9425 438 9535 4 gnd
rlabel metal2 s 330 4939 438 5015 4 gnd
rlabel metal2 s 330 3359 438 3435 4 gnd
rlabel metal2 s 330 9995 438 10071 4 gnd
rlabel metal2 s 330 4685 438 4795 4 gnd
rlabel metal2 s 330 13375 438 13485 4 gnd
rlabel metal2 s 330 10785 438 10861 4 gnd
rlabel metal2 s 330 5255 438 5331 4 gnd
rlabel metal2 s 330 25005 438 25081 4 gnd
rlabel metal2 s 330 16535 438 16645 4 gnd
rlabel metal2 s 330 9679 438 9755 4 gnd
rlabel metal2 s 330 24689 438 24765 4 gnd
rlabel metal2 s 330 13945 438 14021 4 gnd
rlabel metal2 s 330 17895 438 17971 4 gnd
rlabel metal2 s 330 8099 438 8175 4 gnd
rlabel metal2 s 330 4465 438 4541 4 gnd
rlabel metal2 s 330 2315 438 2425 4 gnd
rlabel metal2 s 330 23109 438 23185 4 gnd
rlabel metal2 s 330 6045 438 6121 4 gnd
rlabel metal2 s 330 11259 438 11335 4 gnd
rlabel metal2 s 330 25479 438 25555 4 gnd
rlabel metal2 s 330 11575 438 11651 4 gnd
rlabel metal2 s 330 1305 438 1381 4 gnd
rlabel metal2 s 330 11005 438 11115 4 gnd
rlabel metal2 s 330 19159 438 19235 4 gnd
rlabel metal2 s 330 18369 438 18445 4 gnd
rlabel metal2 s 330 23425 438 23501 4 gnd
rlabel metal2 s 330 14735 438 14811 4 gnd
rlabel metal2 s 330 13155 438 13231 4 gnd
rlabel metal2 s 330 24435 438 24545 4 gnd
rlabel metal2 s 330 18115 438 18225 4 gnd
rlabel metal2 s 330 23899 438 23975 4 gnd
rlabel metal2 s 330 7845 438 7955 4 gnd
rlabel metal2 s 330 3895 438 4005 4 gnd
rlabel metal2 s 330 21529 438 21605 4 gnd
rlabel metal2 s 330 22635 438 22711 4 gnd
rlabel metal2 s 330 16789 438 16865 4 gnd
rlabel metal2 s 330 3105 438 3215 4 gnd
rlabel metal2 s 330 10469 438 10545 4 gnd
rlabel metal2 s 330 16315 438 16391 4 gnd
rlabel metal2 s 330 19695 438 19805 4 gnd
rlabel metal2 s 330 20265 438 20341 4 gnd
rlabel metal2 s 330 25225 438 25335 4 gnd
rlabel metal2 s 330 8635 438 8745 4 gnd
rlabel metal2 s 330 21055 438 21131 4 gnd
rlabel metal2 s 330 6835 438 6911 4 gnd
rlabel metal2 s 330 12585 438 12695 4 gnd
rlabel metal2 s 330 21845 438 21921 4 gnd
rlabel metal2 s 330 5475 438 5585 4 gnd
rlabel metal2 s 330 1779 438 1855 4 gnd
rlabel metal2 s 330 11795 438 11905 4 gnd
rlabel metal2 s 330 17105 438 17181 4 gnd
rlabel metal2 s 330 7309 438 7385 4 gnd
rlabel metal2 s 330 989 438 1065 4 gnd
rlabel metal2 s 330 23645 438 23755 4 gnd
rlabel metal2 s 330 15209 438 15285 4 gnd
rlabel metal2 s 330 18685 438 18761 4 gnd
rlabel metal2 s 330 22319 438 22395 4 gnd
rlabel metal2 s 330 2569 438 2645 4 gnd
rlabel metal2 s 330 4149 438 4225 4 gnd
rlabel metal2 s 330 22065 438 22175 4 gnd
rlabel metal2 s 330 19949 438 20025 4 gnd
rlabel metal2 s 330 17579 438 17655 4 gnd
rlabel metal2 s 330 8889 438 8965 4 gnd
rlabel metal2 s 330 19475 438 19551 4 gnd
rlabel metal2 s 330 735 438 845 4 gnd
rlabel metal2 s 330 6265 438 6375 4 gnd
rlabel metal2 s 330 20739 438 20815 4 gnd
rlabel metal2 s 330 15525 438 15601 4 gnd
rlabel metal2 s 330 12365 438 12441 4 gnd
rlabel metal2 s 330 9205 438 9281 4 gnd
rlabel metal2 s 330 3675 438 3751 4 gnd
rlabel metal2 s 330 14955 438 15065 4 gnd
rlabel metal2 s 330 12839 438 12915 4 gnd
rlabel metal2 s 330 5729 438 5805 4 gnd
rlabel metal2 s 330 22855 438 22965 4 gnd
rlabel metal2 s 330 13629 438 13705 4 gnd
rlabel metal2 s 330 18905 438 19015 4 gnd
rlabel metal2 s 330 1525 438 1635 4 gnd
rlabel metal2 s 330 2885 438 2961 4 gnd
rlabel metal2 s 330 7625 438 7701 4 gnd
rlabel metal2 s 330 2095 438 2171 4 gnd
rlabel metal2 s 330 17325 438 17435 4 gnd
rlabel metal2 s 330 7055 438 7165 4 gnd
rlabel metal2 s 330 20485 438 20595 4 gnd
rlabel metal2 s 330 515 438 591 4 gnd
rlabel metal2 s 330 10215 438 10325 4 gnd
rlabel metal2 s 330 21275 438 21385 4 gnd
rlabel metal2 s 330 24215 438 24291 4 gnd
rlabel metal2 s 330 25795 438 25871 4 gnd
rlabel metal2 s 330 26015 438 26125 4 gnd
rlabel metal2 s 330 8415 438 8491 4 gnd
rlabel metal2 s 330 15745 438 15855 4 gnd
rlabel metal2 s 330 6519 438 6595 4 gnd
rlabel metal2 s 330 14165 438 14275 4 gnd
rlabel metal2 s 330 12049 438 12125 4 gnd
rlabel metal2 s 330 15999 438 16075 4 gnd
rlabel metal2 s 330 14419 438 14495 4 gnd
rlabel metal1 s 366 50639 402 50980 4 vdd
rlabel metal1 s 366 26440 402 26781 4 vdd
rlabel metal1 s 366 28810 402 29151 4 vdd
rlabel metal1 s 366 48560 402 48901 4 vdd
rlabel metal1 s 366 50930 402 51271 4 vdd
rlabel metal1 s 366 29309 402 29650 4 vdd
rlabel metal1 s 366 30889 402 31230 4 vdd
rlabel metal1 s 366 47770 402 48111 4 vdd
rlabel metal1 s 366 43529 402 43870 4 vdd
rlabel metal1 s 366 46689 402 47030 4 vdd
rlabel metal1 s 366 39080 402 39421 4 vdd
rlabel metal1 s 366 43820 402 44161 4 vdd
rlabel metal1 s 366 45400 402 45741 4 vdd
rlabel metal1 s 366 33550 402 33891 4 vdd
rlabel metal1 s 366 34839 402 35180 4 vdd
rlabel metal1 s 366 44610 402 44951 4 vdd
rlabel metal1 s 366 28020 402 28361 4 vdd
rlabel metal1 s 366 44319 402 44660 4 vdd
rlabel metal1 s 366 26149 402 26490 4 vdd
rlabel metal1 s 366 29600 402 29941 4 vdd
rlabel metal1 s 366 36710 402 37051 4 vdd
rlabel metal1 s 366 48269 402 48610 4 vdd
rlabel metal1 s 366 37500 402 37841 4 vdd
rlabel metal1 s 366 41450 402 41791 4 vdd
rlabel metal1 s 366 31970 402 32311 4 vdd
rlabel metal1 s 366 47479 402 47820 4 vdd
rlabel metal1 s 366 51429 402 51770 4 vdd
rlabel metal1 s 366 45899 402 46240 4 vdd
rlabel metal1 s 366 27230 402 27571 4 vdd
rlabel metal1 s 366 37209 402 37550 4 vdd
rlabel metal1 s 366 31679 402 32020 4 vdd
rlabel metal1 s 366 32469 402 32810 4 vdd
rlabel metal1 s 366 38290 402 38631 4 vdd
rlabel metal1 s 366 30390 402 30731 4 vdd
rlabel metal1 s 366 49350 402 49691 4 vdd
rlabel metal1 s 366 26939 402 27280 4 vdd
rlabel metal1 s 366 38789 402 39130 4 vdd
rlabel metal1 s 366 39870 402 40211 4 vdd
rlabel metal1 s 366 49059 402 49400 4 vdd
rlabel metal1 s 366 35130 402 35471 4 vdd
rlabel metal1 s 366 37999 402 38340 4 vdd
rlabel metal1 s 366 41949 402 42290 4 vdd
rlabel metal1 s 366 41159 402 41500 4 vdd
rlabel metal1 s 366 42240 402 42581 4 vdd
rlabel metal1 s 366 46980 402 47321 4 vdd
rlabel metal1 s 366 27729 402 28070 4 vdd
rlabel metal1 s 366 43030 402 43371 4 vdd
rlabel metal1 s 366 46190 402 46531 4 vdd
rlabel metal1 s 366 40660 402 41001 4 vdd
rlabel metal1 s 366 45109 402 45450 4 vdd
rlabel metal1 s 366 36419 402 36760 4 vdd
rlabel metal1 s 366 35920 402 36261 4 vdd
rlabel metal1 s 366 49849 402 50190 4 vdd
rlabel metal1 s 366 42739 402 43080 4 vdd
rlabel metal1 s 366 32760 402 33101 4 vdd
rlabel metal1 s 366 30099 402 30440 4 vdd
rlabel metal1 s 366 35629 402 35970 4 vdd
rlabel metal1 s 366 34049 402 34390 4 vdd
rlabel metal1 s 366 34340 402 34681 4 vdd
rlabel metal1 s 366 39579 402 39920 4 vdd
rlabel metal1 s 366 28519 402 28860 4 vdd
rlabel metal1 s 366 31180 402 31521 4 vdd
rlabel metal1 s 366 40369 402 40710 4 vdd
rlabel metal1 s 366 33259 402 33600 4 vdd
rlabel metal1 s 366 50140 402 50481 4 vdd
rlabel metal1 s 222 0 258 52140 4 br_1_0
rlabel metal1 s 366 18249 402 18590 4 vdd
rlabel metal1 s 366 12719 402 13060 4 vdd
rlabel metal1 s 366 24860 402 25201 4 vdd
rlabel metal1 s 366 7979 402 8320 4 vdd
rlabel metal1 s 366 23779 402 24120 4 vdd
rlabel metal1 s 366 11430 402 11771 4 vdd
rlabel metal1 s 510 0 546 52140 4 bl_0_0
rlabel metal1 s 438 0 474 52140 4 br_0_0
rlabel metal1 s 366 4320 402 4661 4 vdd
rlabel metal1 s 366 22199 402 22540 4 vdd
rlabel metal1 s 366 24569 402 24910 4 vdd
rlabel metal1 s 294 0 330 52140 4 bl_1_0
rlabel metal1 s 366 8769 402 9110 4 vdd
rlabel metal1 s 366 6690 402 7031 4 vdd
rlabel metal1 s 366 13800 402 14141 4 vdd
rlabel metal1 s 366 7189 402 7530 4 vdd
rlabel metal1 s 366 22989 402 23330 4 vdd
rlabel metal1 s 366 4819 402 5160 4 vdd
rlabel metal1 s 366 5110 402 5451 4 vdd
rlabel metal1 s 366 19829 402 20170 4 vdd
rlabel metal1 s 366 3530 402 3871 4 vdd
rlabel metal1 s 366 2449 402 2790 4 vdd
rlabel metal1 s 366 15380 402 15721 4 vdd
rlabel metal1 s 366 21700 402 22041 4 vdd
rlabel metal1 s 366 25359 402 25700 4 vdd
rlabel metal1 s 366 25650 402 25991 4 vdd
rlabel metal1 s 366 16960 402 17301 4 vdd
rlabel metal1 s 366 16170 402 16511 4 vdd
rlabel metal1 s 366 5900 402 6241 4 vdd
rlabel metal1 s 366 20619 402 20960 4 vdd
rlabel metal1 s 366 7480 402 7821 4 vdd
rlabel metal1 s 366 14590 402 14931 4 vdd
rlabel metal1 s 366 11929 402 12270 4 vdd
rlabel metal1 s 366 2740 402 3081 4 vdd
rlabel metal1 s 366 19039 402 19380 4 vdd
rlabel metal1 s 366 20910 402 21251 4 vdd
rlabel metal1 s 366 17459 402 17800 4 vdd
rlabel metal1 s 366 15879 402 16220 4 vdd
rlabel metal1 s 366 1659 402 2000 4 vdd
rlabel metal1 s 366 4029 402 4370 4 vdd
rlabel metal1 s 366 13010 402 13351 4 vdd
rlabel metal1 s 366 24070 402 24411 4 vdd
rlabel metal1 s 366 17750 402 18091 4 vdd
rlabel metal1 s 366 22490 402 22831 4 vdd
rlabel metal1 s 366 9850 402 10191 4 vdd
rlabel metal1 s 366 16669 402 17010 4 vdd
rlabel metal1 s 366 20120 402 20461 4 vdd
rlabel metal1 s 366 9060 402 9401 4 vdd
rlabel metal1 s 366 370 402 711 4 vdd
rlabel metal1 s 366 3239 402 3580 4 vdd
rlabel metal1 s 366 19330 402 19671 4 vdd
rlabel metal1 s 366 1160 402 1501 4 vdd
rlabel metal1 s 366 15089 402 15430 4 vdd
rlabel metal1 s 366 13509 402 13850 4 vdd
rlabel metal1 s 366 869 402 1210 4 vdd
rlabel metal1 s 366 10349 402 10690 4 vdd
rlabel metal1 s 366 1950 402 2291 4 vdd
rlabel metal1 s 366 21409 402 21750 4 vdd
rlabel metal1 s 366 8270 402 8611 4 vdd
rlabel metal1 s 366 10640 402 10981 4 vdd
rlabel metal1 s 366 5609 402 5950 4 vdd
rlabel metal1 s 366 23280 402 23621 4 vdd
rlabel metal1 s 366 9559 402 9900 4 vdd
rlabel metal1 s 366 11139 402 11480 4 vdd
rlabel metal1 s 366 6399 402 6740 4 vdd
rlabel metal1 s 366 18540 402 18881 4 vdd
rlabel metal1 s 366 14299 402 14640 4 vdd
rlabel metal1 s 366 12220 402 12561 4 vdd
<< properties >>
string FIXED_BBOX 0 0 624 52140
string GDS_END 1799030
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 1683822
<< end >>
