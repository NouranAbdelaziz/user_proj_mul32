/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/klayout/pymacros/cells/fixed_devices/VPP/sky130_fd_pr__cap_vpp_11p5x11p7_m1m4_noshield.cdl