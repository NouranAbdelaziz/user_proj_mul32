magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< pwell >>
rect 10 10 634 662
<< nmoslvt >>
rect 92 36 122 636
rect 178 36 208 636
rect 264 36 294 636
rect 350 36 380 636
rect 436 36 466 636
rect 522 36 552 636
<< ndiff >>
rect 36 605 92 636
rect 36 571 47 605
rect 81 571 92 605
rect 36 533 92 571
rect 36 499 47 533
rect 81 499 92 533
rect 36 461 92 499
rect 36 427 47 461
rect 81 427 92 461
rect 36 389 92 427
rect 36 355 47 389
rect 81 355 92 389
rect 36 317 92 355
rect 36 283 47 317
rect 81 283 92 317
rect 36 245 92 283
rect 36 211 47 245
rect 81 211 92 245
rect 36 173 92 211
rect 36 139 47 173
rect 81 139 92 173
rect 36 101 92 139
rect 36 67 47 101
rect 81 67 92 101
rect 36 36 92 67
rect 122 605 178 636
rect 122 571 133 605
rect 167 571 178 605
rect 122 533 178 571
rect 122 499 133 533
rect 167 499 178 533
rect 122 461 178 499
rect 122 427 133 461
rect 167 427 178 461
rect 122 389 178 427
rect 122 355 133 389
rect 167 355 178 389
rect 122 317 178 355
rect 122 283 133 317
rect 167 283 178 317
rect 122 245 178 283
rect 122 211 133 245
rect 167 211 178 245
rect 122 173 178 211
rect 122 139 133 173
rect 167 139 178 173
rect 122 101 178 139
rect 122 67 133 101
rect 167 67 178 101
rect 122 36 178 67
rect 208 605 264 636
rect 208 571 219 605
rect 253 571 264 605
rect 208 533 264 571
rect 208 499 219 533
rect 253 499 264 533
rect 208 461 264 499
rect 208 427 219 461
rect 253 427 264 461
rect 208 389 264 427
rect 208 355 219 389
rect 253 355 264 389
rect 208 317 264 355
rect 208 283 219 317
rect 253 283 264 317
rect 208 245 264 283
rect 208 211 219 245
rect 253 211 264 245
rect 208 173 264 211
rect 208 139 219 173
rect 253 139 264 173
rect 208 101 264 139
rect 208 67 219 101
rect 253 67 264 101
rect 208 36 264 67
rect 294 605 350 636
rect 294 571 305 605
rect 339 571 350 605
rect 294 533 350 571
rect 294 499 305 533
rect 339 499 350 533
rect 294 461 350 499
rect 294 427 305 461
rect 339 427 350 461
rect 294 389 350 427
rect 294 355 305 389
rect 339 355 350 389
rect 294 317 350 355
rect 294 283 305 317
rect 339 283 350 317
rect 294 245 350 283
rect 294 211 305 245
rect 339 211 350 245
rect 294 173 350 211
rect 294 139 305 173
rect 339 139 350 173
rect 294 101 350 139
rect 294 67 305 101
rect 339 67 350 101
rect 294 36 350 67
rect 380 605 436 636
rect 380 571 391 605
rect 425 571 436 605
rect 380 533 436 571
rect 380 499 391 533
rect 425 499 436 533
rect 380 461 436 499
rect 380 427 391 461
rect 425 427 436 461
rect 380 389 436 427
rect 380 355 391 389
rect 425 355 436 389
rect 380 317 436 355
rect 380 283 391 317
rect 425 283 436 317
rect 380 245 436 283
rect 380 211 391 245
rect 425 211 436 245
rect 380 173 436 211
rect 380 139 391 173
rect 425 139 436 173
rect 380 101 436 139
rect 380 67 391 101
rect 425 67 436 101
rect 380 36 436 67
rect 466 605 522 636
rect 466 571 477 605
rect 511 571 522 605
rect 466 533 522 571
rect 466 499 477 533
rect 511 499 522 533
rect 466 461 522 499
rect 466 427 477 461
rect 511 427 522 461
rect 466 389 522 427
rect 466 355 477 389
rect 511 355 522 389
rect 466 317 522 355
rect 466 283 477 317
rect 511 283 522 317
rect 466 245 522 283
rect 466 211 477 245
rect 511 211 522 245
rect 466 173 522 211
rect 466 139 477 173
rect 511 139 522 173
rect 466 101 522 139
rect 466 67 477 101
rect 511 67 522 101
rect 466 36 522 67
rect 552 605 608 636
rect 552 571 563 605
rect 597 571 608 605
rect 552 533 608 571
rect 552 499 563 533
rect 597 499 608 533
rect 552 461 608 499
rect 552 427 563 461
rect 597 427 608 461
rect 552 389 608 427
rect 552 355 563 389
rect 597 355 608 389
rect 552 317 608 355
rect 552 283 563 317
rect 597 283 608 317
rect 552 245 608 283
rect 552 211 563 245
rect 597 211 608 245
rect 552 173 608 211
rect 552 139 563 173
rect 597 139 608 173
rect 552 101 608 139
rect 552 67 563 101
rect 597 67 608 101
rect 552 36 608 67
<< ndiffc >>
rect 47 571 81 605
rect 47 499 81 533
rect 47 427 81 461
rect 47 355 81 389
rect 47 283 81 317
rect 47 211 81 245
rect 47 139 81 173
rect 47 67 81 101
rect 133 571 167 605
rect 133 499 167 533
rect 133 427 167 461
rect 133 355 167 389
rect 133 283 167 317
rect 133 211 167 245
rect 133 139 167 173
rect 133 67 167 101
rect 219 571 253 605
rect 219 499 253 533
rect 219 427 253 461
rect 219 355 253 389
rect 219 283 253 317
rect 219 211 253 245
rect 219 139 253 173
rect 219 67 253 101
rect 305 571 339 605
rect 305 499 339 533
rect 305 427 339 461
rect 305 355 339 389
rect 305 283 339 317
rect 305 211 339 245
rect 305 139 339 173
rect 305 67 339 101
rect 391 571 425 605
rect 391 499 425 533
rect 391 427 425 461
rect 391 355 425 389
rect 391 283 425 317
rect 391 211 425 245
rect 391 139 425 173
rect 391 67 425 101
rect 477 571 511 605
rect 477 499 511 533
rect 477 427 511 461
rect 477 355 511 389
rect 477 283 511 317
rect 477 211 511 245
rect 477 139 511 173
rect 477 67 511 101
rect 563 571 597 605
rect 563 499 597 533
rect 563 427 597 461
rect 563 355 597 389
rect 563 283 597 317
rect 563 211 597 245
rect 563 139 597 173
rect 563 67 597 101
<< poly >>
rect 92 717 552 733
rect 92 683 135 717
rect 169 683 203 717
rect 237 683 271 717
rect 305 683 339 717
rect 373 683 407 717
rect 441 683 475 717
rect 509 683 552 717
rect 92 662 552 683
rect 92 636 122 662
rect 178 636 208 662
rect 264 636 294 662
rect 350 636 380 662
rect 436 636 466 662
rect 522 636 552 662
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
rect 436 10 466 36
rect 522 10 552 36
<< polycont >>
rect 135 683 169 717
rect 203 683 237 717
rect 271 683 305 717
rect 339 683 373 717
rect 407 683 441 717
rect 475 683 509 717
<< locali >>
rect 119 717 525 733
rect 119 683 125 717
rect 169 683 197 717
rect 237 683 269 717
rect 305 683 339 717
rect 375 683 407 717
rect 447 683 475 717
rect 519 683 525 717
rect 119 667 525 683
rect 47 605 81 621
rect 47 533 81 571
rect 47 461 81 499
rect 47 389 81 427
rect 47 317 81 355
rect 47 245 81 283
rect 47 173 81 211
rect 47 101 81 139
rect 47 51 81 67
rect 133 605 167 621
rect 133 533 167 571
rect 133 461 167 499
rect 133 389 167 427
rect 133 317 167 355
rect 133 245 167 283
rect 133 173 167 211
rect 133 101 167 139
rect 133 51 167 67
rect 219 605 253 621
rect 219 533 253 571
rect 219 461 253 499
rect 219 389 253 427
rect 219 317 253 355
rect 219 245 253 283
rect 219 173 253 211
rect 219 101 253 139
rect 219 51 253 67
rect 305 605 339 621
rect 305 533 339 571
rect 305 461 339 499
rect 305 389 339 427
rect 305 317 339 355
rect 305 245 339 283
rect 305 173 339 211
rect 305 101 339 139
rect 305 51 339 67
rect 391 605 425 621
rect 391 533 425 571
rect 391 461 425 499
rect 391 389 425 427
rect 391 317 425 355
rect 391 245 425 283
rect 391 173 425 211
rect 391 101 425 139
rect 391 51 425 67
rect 477 605 511 621
rect 477 533 511 571
rect 477 461 511 499
rect 477 389 511 427
rect 477 317 511 355
rect 477 245 511 283
rect 477 173 511 211
rect 477 101 511 139
rect 477 51 511 67
rect 563 605 597 621
rect 563 533 597 571
rect 563 461 597 499
rect 563 389 597 427
rect 563 317 597 355
rect 563 245 597 283
rect 563 173 597 211
rect 563 101 597 139
rect 563 51 597 67
<< viali >>
rect 125 683 135 717
rect 135 683 159 717
rect 197 683 203 717
rect 203 683 231 717
rect 269 683 271 717
rect 271 683 303 717
rect 341 683 373 717
rect 373 683 375 717
rect 413 683 441 717
rect 441 683 447 717
rect 485 683 509 717
rect 509 683 519 717
rect 47 571 81 605
rect 47 499 81 533
rect 47 427 81 461
rect 47 355 81 389
rect 47 283 81 317
rect 47 211 81 245
rect 47 139 81 173
rect 47 67 81 101
rect 133 571 167 605
rect 133 499 167 533
rect 133 427 167 461
rect 133 355 167 389
rect 133 283 167 317
rect 133 211 167 245
rect 133 139 167 173
rect 133 67 167 101
rect 219 571 253 605
rect 219 499 253 533
rect 219 427 253 461
rect 219 355 253 389
rect 219 283 253 317
rect 219 211 253 245
rect 219 139 253 173
rect 219 67 253 101
rect 305 571 339 605
rect 305 499 339 533
rect 305 427 339 461
rect 305 355 339 389
rect 305 283 339 317
rect 305 211 339 245
rect 305 139 339 173
rect 305 67 339 101
rect 391 571 425 605
rect 391 499 425 533
rect 391 427 425 461
rect 391 355 425 389
rect 391 283 425 317
rect 391 211 425 245
rect 391 139 425 173
rect 391 67 425 101
rect 477 571 511 605
rect 477 499 511 533
rect 477 427 511 461
rect 477 355 511 389
rect 477 283 511 317
rect 477 211 511 245
rect 477 139 511 173
rect 477 67 511 101
rect 563 571 597 605
rect 563 499 597 533
rect 563 427 597 461
rect 563 355 597 389
rect 563 283 597 317
rect 563 211 597 245
rect 563 139 597 173
rect 563 67 597 101
<< metal1 >>
rect 113 717 531 729
rect 113 683 125 717
rect 159 683 197 717
rect 231 683 269 717
rect 303 683 341 717
rect 375 683 413 717
rect 447 683 485 717
rect 519 683 531 717
rect 113 671 531 683
rect 41 605 87 621
rect 41 571 47 605
rect 81 571 87 605
rect 41 533 87 571
rect 41 499 47 533
rect 81 499 87 533
rect 41 461 87 499
rect 41 427 47 461
rect 81 427 87 461
rect 41 389 87 427
rect 41 355 47 389
rect 81 355 87 389
rect 41 317 87 355
rect 41 283 47 317
rect 81 283 87 317
rect 41 245 87 283
rect 41 211 47 245
rect 81 211 87 245
rect 41 173 87 211
rect 41 139 47 173
rect 81 139 87 173
rect 41 101 87 139
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 124 608 176 621
rect 124 544 176 556
rect 124 461 176 492
rect 124 427 133 461
rect 167 427 176 461
rect 124 389 176 427
rect 124 355 133 389
rect 167 355 176 389
rect 124 317 176 355
rect 124 283 133 317
rect 167 283 176 317
rect 124 245 176 283
rect 124 211 133 245
rect 167 211 176 245
rect 124 173 176 211
rect 124 139 133 173
rect 167 139 176 173
rect 124 101 176 139
rect 124 67 133 101
rect 167 67 176 101
rect 124 51 176 67
rect 213 605 259 621
rect 213 571 219 605
rect 253 571 259 605
rect 213 533 259 571
rect 213 499 219 533
rect 253 499 259 533
rect 213 461 259 499
rect 213 427 219 461
rect 253 427 259 461
rect 213 389 259 427
rect 213 355 219 389
rect 253 355 259 389
rect 213 317 259 355
rect 213 283 219 317
rect 253 283 259 317
rect 213 245 259 283
rect 213 211 219 245
rect 253 211 259 245
rect 213 173 259 211
rect 213 139 219 173
rect 253 139 259 173
rect 213 101 259 139
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 296 608 348 621
rect 296 544 348 556
rect 296 461 348 492
rect 296 427 305 461
rect 339 427 348 461
rect 296 389 348 427
rect 296 355 305 389
rect 339 355 348 389
rect 296 317 348 355
rect 296 283 305 317
rect 339 283 348 317
rect 296 245 348 283
rect 296 211 305 245
rect 339 211 348 245
rect 296 173 348 211
rect 296 139 305 173
rect 339 139 348 173
rect 296 101 348 139
rect 296 67 305 101
rect 339 67 348 101
rect 296 51 348 67
rect 385 605 431 621
rect 385 571 391 605
rect 425 571 431 605
rect 385 533 431 571
rect 385 499 391 533
rect 425 499 431 533
rect 385 461 431 499
rect 385 427 391 461
rect 425 427 431 461
rect 385 389 431 427
rect 385 355 391 389
rect 425 355 431 389
rect 385 317 431 355
rect 385 283 391 317
rect 425 283 431 317
rect 385 245 431 283
rect 385 211 391 245
rect 425 211 431 245
rect 385 173 431 211
rect 385 139 391 173
rect 425 139 431 173
rect 385 101 431 139
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 468 608 520 621
rect 468 544 520 556
rect 468 461 520 492
rect 468 427 477 461
rect 511 427 520 461
rect 468 389 520 427
rect 468 355 477 389
rect 511 355 520 389
rect 468 317 520 355
rect 468 283 477 317
rect 511 283 520 317
rect 468 245 520 283
rect 468 211 477 245
rect 511 211 520 245
rect 468 173 520 211
rect 468 139 477 173
rect 511 139 520 173
rect 468 101 520 139
rect 468 67 477 101
rect 511 67 520 101
rect 468 51 520 67
rect 557 605 603 621
rect 557 571 563 605
rect 597 571 603 605
rect 557 533 603 571
rect 557 499 563 533
rect 597 499 603 533
rect 557 461 603 499
rect 557 427 563 461
rect 597 427 603 461
rect 557 389 603 427
rect 557 355 563 389
rect 597 355 603 389
rect 557 317 603 355
rect 557 283 563 317
rect 597 283 603 317
rect 557 245 603 283
rect 557 211 563 245
rect 597 211 603 245
rect 557 173 603 211
rect 557 139 563 173
rect 597 139 603 173
rect 557 101 603 139
rect 557 67 563 101
rect 597 67 603 101
rect 557 -29 603 67
rect 41 -89 603 -29
<< via1 >>
rect 124 605 176 608
rect 124 571 133 605
rect 133 571 167 605
rect 167 571 176 605
rect 124 556 176 571
rect 124 533 176 544
rect 124 499 133 533
rect 133 499 167 533
rect 167 499 176 533
rect 124 492 176 499
rect 296 605 348 608
rect 296 571 305 605
rect 305 571 339 605
rect 339 571 348 605
rect 296 556 348 571
rect 296 533 348 544
rect 296 499 305 533
rect 305 499 339 533
rect 339 499 348 533
rect 296 492 348 499
rect 468 605 520 608
rect 468 571 477 605
rect 477 571 511 605
rect 511 571 520 605
rect 468 556 520 571
rect 468 533 520 544
rect 468 499 477 533
rect 477 499 511 533
rect 511 499 520 533
rect 468 492 520 499
<< metal2 >>
rect 117 618 183 627
rect 117 562 122 618
rect 178 562 183 618
rect 117 556 124 562
rect 176 556 183 562
rect 117 544 183 556
rect 117 538 124 544
rect 176 538 183 544
rect 117 482 122 538
rect 178 482 183 538
rect 117 473 183 482
rect 289 618 355 627
rect 289 562 294 618
rect 350 562 355 618
rect 289 556 296 562
rect 348 556 355 562
rect 289 544 355 556
rect 289 538 296 544
rect 348 538 355 544
rect 289 482 294 538
rect 350 482 355 538
rect 289 473 355 482
rect 461 618 527 627
rect 461 562 466 618
rect 522 562 527 618
rect 461 556 468 562
rect 520 556 527 562
rect 461 544 527 556
rect 461 538 468 544
rect 520 538 527 544
rect 461 482 466 538
rect 522 482 527 538
rect 461 473 527 482
<< via2 >>
rect 122 608 178 618
rect 122 562 124 608
rect 124 562 176 608
rect 176 562 178 608
rect 122 492 124 538
rect 124 492 176 538
rect 176 492 178 538
rect 122 482 178 492
rect 294 608 350 618
rect 294 562 296 608
rect 296 562 348 608
rect 348 562 350 608
rect 294 492 296 538
rect 296 492 348 538
rect 348 492 350 538
rect 294 482 350 492
rect 466 608 522 618
rect 466 562 468 608
rect 468 562 520 608
rect 520 562 522 608
rect 466 492 468 538
rect 468 492 520 538
rect 520 492 522 538
rect 466 482 522 492
<< metal3 >>
rect 117 618 527 627
rect 117 562 122 618
rect 178 562 294 618
rect 350 562 466 618
rect 522 562 527 618
rect 117 561 527 562
rect 117 538 183 561
rect 117 482 122 538
rect 178 482 183 538
rect 117 473 183 482
rect 289 538 355 561
rect 289 482 294 538
rect 350 482 355 538
rect 289 473 355 482
rect 461 538 527 561
rect 461 482 466 538
rect 522 482 527 538
rect 461 473 527 482
<< labels >>
flabel metal3 s 117 561 527 627 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 41 -89 603 -29 0 FreeSans 400 0 0 0 SOURCE
port 2 nsew
flabel metal1 s 113 671 531 729 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel pwell s 72 641 90 653 0 FreeSans 200 0 0 0 SUBSTRATE
<< properties >>
string GDS_END 3374310
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3359464
string path 1.600 15.525 1.600 -2.225 
<< end >>
