/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/parasitics/sky130_fd_pr__model__parasitic__diode_pw2dn__extended_drain.model.spice