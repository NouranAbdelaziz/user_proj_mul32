/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/klayout/pymacros/cells/fixed_devices/VPP/sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x8.cdl