magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< obsactive >>
tri 25423 26223 40000 40800 ne
<< metal4 >>
rect 0 35957 254 40800
rect 0 14807 254 19800
rect 0 13617 254 14507
rect 0 12447 254 13337
rect 0 12081 254 12147
rect 0 11425 100 12021
rect 0 11129 254 11365
rect 0 10473 116 11069
rect 0 10347 254 10413
rect 0 9117 254 10047
rect 0 8147 254 8837
rect 0 7177 254 7867
rect 0 5967 254 6897
rect 0 4757 254 5687
rect 0 3787 254 4477
rect 0 2577 254 3507
rect 0 1207 254 2297
rect 407 0 1497 254
rect 1777 0 2707 254
rect 2987 0 3677 254
rect 3957 0 4887 254
rect 5167 0 6097 254
rect 6377 0 7067 254
rect 7347 0 8037 254
rect 8317 0 9247 254
rect 9547 0 9613 254
rect 9673 0 10269 115
rect 10329 0 10565 254
rect 10625 0 11221 100
rect 11281 0 11347 254
rect 11647 0 12537 254
rect 12817 0 13707 254
rect 14007 0 19000 254
rect 35157 0 40000 254
<< metal5 >>
rect 0 35957 254 40800
rect 0 14807 254 19797
rect 0 13637 254 14487
rect 0 12467 254 13317
rect 0 10347 254 12147
rect 0 9137 254 10027
rect 0 8167 254 8817
rect 0 7197 254 7847
rect 0 5987 254 6877
rect 0 4777 254 5667
rect 0 3807 254 4457
rect 0 2597 254 3487
rect 0 1227 254 2277
rect 427 0 1477 254
rect 1797 0 2687 254
rect 3007 0 3657 254
rect 3977 0 4867 254
rect 5187 0 6077 254
rect 6397 0 7047 254
rect 7367 0 8017 254
rect 8337 0 9227 254
rect 9547 0 11347 254
rect 11667 0 12517 254
rect 12837 0 13687 254
rect 14007 0 18997 254
rect 35157 0 40000 254
<< fillblock >>
tri 25423 26223 40000 40800 ne
use sky130_fd_io__corner_bus_overlay  sky130_fd_io__corner_bus_overlay_0
timestamp 1676037725
transform 1 0 0 0 1 67
box 0 0 40000 40733
<< labels >>
flabel metal4 s 0 11425 100 12021 3 FreeSans 650 0 0 0 AMUXBUS_A
flabel metal4 s 10625 0 11221 100 3 FreeSans 650 90 0 0 AMUXBUS_A
port 1 e
flabel metal4 s 0 10473 115 11069 3 FreeSans 650 0 0 0 AMUXBUS_B
flabel metal4 s 9673 0 10269 115 3 FreeSans 650 90 0 0 AMUXBUS_B
port 2 e
flabel metal5 s 0 10347 254 12147 3 FreeSans 650 0 0 0 VSSA
flabel metal5 s 127 11205 127 11205 3 FreeSans 650 180 0 0 VSSA
flabel metal5 s 0 8168 254 8817 3 FreeSans 650 180 0 0 VSSA
flabel metal4 s 0 10347 254 10413 3 FreeSans 650 0 0 0 VSSA
flabel metal4 s 0 8147 254 8837 3 FreeSans 650 180 0 0 VSSA
flabel metal4 s 0 11129 254 11365 3 FreeSans 650 0 0 0 VSSA
flabel metal4 s 0 12081 254 12147 3 FreeSans 650 0 0 0 VSSA
flabel metal5 s 7368 0 8017 254 3 FreeSans 650 270 0 0 VSSA
flabel metal5 s 9547 0 11347 254 3 FreeSans 650 270 0 0 VSSA
flabel metal5 s 10258 127 10258 127 3 FreeSans 650 90 0 0 VSSA
flabel metal4 s 11281 0 11347 254 3 FreeSans 650 90 0 0 VSSA
flabel metal4 s 10329 0 10565 254 3 FreeSans 650 90 0 0 VSSA
flabel metal4 s 7347 0 8037 254 3 FreeSans 650 270 0 0 VSSA
flabel metal4 s 9547 0 9613 254 3 FreeSans 650 90 0 0 VSSA
port 3 e
flabel metal5 s 0 3807 251 4457 3 FreeSans 650 180 0 0 VDDA
flabel metal4 s 0 3787 251 4477 3 FreeSans 650 180 0 0 VDDA
flabel metal5 s 3007 0 3657 251 3 FreeSans 650 270 0 0 VDDA
flabel metal4 s 2987 0 3677 251 3 FreeSans 650 270 0 0 VDDA
port 4 e
flabel metal5 s 0 7197 254 7847 3 FreeSans 650 180 0 0 VSWITCH
flabel metal4 s 0 7177 254 7867 3 FreeSans 650 180 0 0 VSWITCH
flabel metal5 s 6397 0 7047 254 3 FreeSans 650 270 0 0 VSWITCH
flabel metal4 s 6377 0 7067 254 3 FreeSans 650 270 0 0 VSWITCH
port 5 e
flabel metal5 s 0 13637 254 14487 3 FreeSans 650 180 0 0 VDDIO_Q
flabel metal4 s 0 13617 254 14507 3 FreeSans 650 180 0 0 VDDIO_Q
flabel metal5 s 12837 0 13687 254 3 FreeSans 650 270 0 0 VDDIO_Q
flabel metal4 s 12817 0 13707 254 3 FreeSans 650 270 0 0 VDDIO_Q
port 6 e
flabel metal5 s 0 1227 254 2277 3 FreeSans 650 180 0 0 VCCHIB
flabel metal4 s 0 1207 254 2297 3 FreeSans 650 180 0 0 VCCHIB
flabel metal5 s 427 0 1477 254 3 FreeSans 650 270 0 0 VCCHIB
flabel metal4 s 407 0 1497 254 3 FreeSans 650 270 0 0 VCCHIB
port 7 e
flabel metal5 s 0 14807 254 19797 3 FreeSans 650 180 0 0 VDDIO
flabel metal5 s 0 4777 254 5667 3 FreeSans 650 180 0 0 VDDIO
flabel metal4 s 0 4757 254 5687 3 FreeSans 650 180 0 0 VDDIO
flabel metal4 s 0 14808 254 19800 3 FreeSans 650 180 0 0 VDDIO
flabel metal5 s 3977 0 4867 254 3 FreeSans 650 270 0 0 VDDIO
flabel metal5 s 14007 0 18997 254 3 FreeSans 650 270 0 0 VDDIO
flabel metal4 s 14008 0 19000 254 3 FreeSans 650 270 0 0 VDDIO
flabel metal4 s 3957 0 4887 254 3 FreeSans 650 270 0 0 VDDIO
port 8 e
flabel metal5 s 0 2597 254 3487 3 FreeSans 650 180 0 0 VCCD
flabel metal4 s 0 2577 254 3507 3 FreeSans 650 180 0 0 VCCD
flabel metal5 s 1797 0 2687 254 3 FreeSans 650 270 0 0 VCCD
flabel metal4 s 1777 0 2707 254 3 FreeSans 650 270 0 0 VCCD
port 9 e
flabel metal5 s 0 5987 254 6877 3 FreeSans 650 180 0 0 VSSIO
flabel metal4 s 0 5967 254 6897 3 FreeSans 650 180 0 0 VSSIO
flabel metal4 s 0 35957 254 40800 3 FreeSans 650 180 0 0 VSSIO
flabel metal4 s 127 38974 127 38974 3 FreeSans 650 180 0 0 VSSIO
flabel metal5 s 5187 0 6077 254 3 FreeSans 650 270 0 0 VSSIO
flabel metal4 s 5167 0 6097 254 3 FreeSans 650 270 0 0 VSSIO
flabel metal4 s 35157 0 40000 254 3 FreeSans 650 270 0 0 VSSIO
flabel metal4 s 38174 127 38174 127 3 FreeSans 650 270 0 0 VSSIO
port 10 e
flabel metal5 s 0 9137 254 10027 3 FreeSans 650 180 0 0 VSSD
flabel metal4 s 0 9117 254 10047 3 FreeSans 650 180 0 0 VSSD
flabel metal5 s 8337 0 9227 254 3 FreeSans 650 270 0 0 VSSD
flabel metal4 s 8317 0 9247 254 3 FreeSans 650 270 0 0 VSSD
port 11 e
flabel metal5 s 0 12467 254 13317 3 FreeSans 650 180 0 0 VSSIO_Q
flabel metal4 s 0 12447 254 13337 3 FreeSans 650 180 0 0 VSSIO_Q
flabel metal5 s 11667 0 12517 254 3 FreeSans 650 270 0 0 VSSIO_Q
flabel metal4 s 11647 0 12537 254 3 FreeSans 650 270 0 0 VSSIO_Q
port 12 e
<< properties >>
string FIXED_BBOX 0 0 40000 40800
string GDS_END 2438082
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 2425268
<< end >>
