/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/sonos_e/end_of_life/typical/ss.spice