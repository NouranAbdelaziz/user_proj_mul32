magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -66 377 1986 897
<< pwell >>
rect 23 43 1901 317
rect -26 -43 1946 43
<< locali >>
rect 127 316 449 363
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 123 729 1901 759
rect 49 453 87 709
rect 157 695 195 729
rect 229 695 267 729
rect 301 695 339 729
rect 373 725 554 729
rect 123 489 373 695
rect 553 695 554 725
rect 588 695 626 729
rect 660 725 821 729
rect 660 695 687 725
rect 409 453 519 689
rect 553 477 687 695
rect 855 695 893 729
rect 927 695 965 729
rect 999 725 1133 729
rect 49 419 519 453
rect 49 295 87 419
rect 485 391 519 419
rect 721 441 787 689
rect 821 477 999 695
rect 1167 695 1205 729
rect 1239 695 1277 729
rect 1311 725 1446 729
rect 1033 441 1099 689
rect 1133 477 1311 695
rect 1445 695 1446 725
rect 1480 695 1589 729
rect 1623 725 1853 729
rect 1781 695 1853 725
rect 1887 695 1901 729
rect 1345 441 1411 689
rect 1445 477 1623 695
rect 1657 646 1747 689
rect 1657 441 1793 646
rect 1827 477 1901 695
rect 721 407 1793 441
rect 485 325 676 391
rect 733 325 1711 359
rect 49 161 91 295
rect 485 280 519 325
rect 135 110 385 277
rect 421 246 519 280
rect 421 146 463 246
rect 553 152 699 289
rect 733 161 775 325
rect 521 110 699 152
rect 809 110 1011 289
rect 1045 161 1087 325
rect 1121 110 1323 289
rect 1357 161 1399 325
rect 1433 110 1635 289
rect 1669 195 1711 325
rect 1747 195 1793 407
rect 1669 161 1793 195
rect 1827 120 1901 289
rect 1795 110 1901 120
rect 135 76 207 110
rect 241 76 279 110
rect 313 76 351 110
rect 385 76 521 110
rect 555 76 593 110
rect 627 76 665 110
rect 699 76 814 110
rect 848 76 886 110
rect 920 76 958 110
rect 992 76 1134 110
rect 1168 76 1206 110
rect 1240 76 1278 110
rect 1312 76 1447 110
rect 1481 76 1519 110
rect 1553 76 1591 110
rect 1625 76 1795 110
rect 1829 76 1867 110
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 123 695 157 729
rect 195 695 229 729
rect 267 695 301 729
rect 339 695 373 729
rect 554 695 588 729
rect 626 695 660 729
rect 821 695 855 729
rect 893 695 927 729
rect 965 695 999 729
rect 1133 695 1167 729
rect 1205 695 1239 729
rect 1277 695 1311 729
rect 1446 695 1480 729
rect 1589 695 1623 729
rect 1853 695 1887 729
rect 207 76 241 110
rect 279 76 313 110
rect 351 76 385 110
rect 521 76 555 110
rect 593 76 627 110
rect 665 76 699 110
rect 814 76 848 110
rect 886 76 920 110
rect 958 76 992 110
rect 1134 76 1168 110
rect 1206 76 1240 110
rect 1278 76 1312 110
rect 1447 76 1481 110
rect 1519 76 1553 110
rect 1591 76 1625 110
rect 1795 76 1829 110
rect 1867 76 1901 110
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 831 1920 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 0 791 1920 797
rect 0 729 1920 763
rect 0 695 123 729
rect 157 695 195 729
rect 229 695 267 729
rect 301 695 339 729
rect 373 695 554 729
rect 588 695 626 729
rect 660 695 821 729
rect 855 695 893 729
rect 927 695 965 729
rect 999 695 1133 729
rect 1167 695 1205 729
rect 1239 695 1277 729
rect 1311 695 1446 729
rect 1480 695 1589 729
rect 1623 695 1853 729
rect 1887 695 1920 729
rect 0 689 1920 695
rect 0 110 1920 125
rect 0 76 207 110
rect 241 76 279 110
rect 313 76 351 110
rect 385 76 521 110
rect 555 76 593 110
rect 627 76 665 110
rect 699 76 814 110
rect 848 76 886 110
rect 920 76 958 110
rect 992 76 1134 110
rect 1168 76 1206 110
rect 1240 76 1278 110
rect 1312 76 1447 110
rect 1481 76 1519 110
rect 1553 76 1591 110
rect 1625 76 1795 110
rect 1829 76 1867 110
rect 1901 76 1920 110
rect 0 51 1920 76
rect 0 17 1920 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -23 1920 -17
<< obsm1 >>
rect 1101 401 1463 447
rect 1101 395 1229 401
<< obsm2 >>
rect 1097 373 1233 447
<< obsm3 >>
rect 1087 377 1243 443
<< obsm4 >>
rect 682 271 1238 507
<< metal5 >>
rect 658 247 1262 567
<< labels >>
rlabel locali s 127 316 449 363 6 A
port 1 nsew signal input
rlabel metal1 s 0 51 1920 125 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 1920 23 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s -26 -43 1946 43 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 23 43 1901 317 6 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 1920 837 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 1986 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 1920 763 6 VPWR
port 5 nsew power bidirectional
rlabel metal5 s 658 247 1262 567 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1920 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 357168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 336410
<< end >>
