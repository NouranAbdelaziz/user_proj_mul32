magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -103 33703 15124 34042
rect -103 29338 335 33703
rect 14619 29338 15124 33703
rect -103 28976 15124 29338
rect -66 26133 15066 28076
<< pwell >>
rect -58 28137 15058 28913
rect -26 25863 8350 26071
rect 12382 25863 15026 26071
rect -26 24827 15026 25863
rect -26 20505 287 24827
rect 14712 20505 15026 24827
rect -26 19846 15026 20505
rect -26 19599 11694 19846
rect 14386 19599 15026 19846
rect -26 19347 15026 19599
rect -26 19346 11694 19347
<< obsli1 >>
rect 0 28887 15000 39844
rect -32 28163 15032 28887
rect 0 26045 15000 28163
rect -53 20279 15000 26045
rect 0 37 15000 20279
<< metal1 >>
rect 2457 0 2509 66
rect 2911 0 3027 66
rect 4472 0 4532 66
rect 4981 0 5027 1995
rect 5516 0 5646 66
rect 6101 0 6231 66
rect 6552 0 6604 66
<< obsm1 >>
rect 0 34018 15000 39842
rect -29 26255 15029 34018
rect 0 26044 15000 26255
rect -29 19179 15029 26044
rect 0 2051 15000 19179
rect 0 122 4925 2051
rect 0 37 2401 122
rect 2565 37 2855 122
rect 3083 37 4416 122
rect 4588 37 4925 122
rect 5083 122 15000 2051
rect 5083 37 5460 122
rect 5702 37 6045 122
rect 6287 37 6496 122
rect 6660 37 15000 122
<< metal2 >>
rect 5864 1072 5916 2217
rect 1685 0 1779 66
rect 2457 0 2509 66
rect 2911 0 3027 66
rect 3449 0 3782 113
rect 4015 0 4245 282
rect 4472 0 4532 66
rect 5516 0 5646 66
rect 5787 0 5933 66
rect 6101 0 6231 66
rect 6552 0 6604 66
rect 14443 0 14647 66
<< obsm2 >>
rect 68 2273 14983 39842
rect 68 1016 5808 2273
rect 5972 1016 14983 2273
rect 68 338 14983 1016
rect 68 169 3959 338
rect 68 122 3393 169
rect 68 0 1629 122
rect 1835 0 2401 122
rect 2565 0 2855 122
rect 3083 0 3393 122
rect 3838 0 3959 169
rect 4301 122 14983 338
rect 4301 0 4416 122
rect 4588 0 5460 122
rect 5702 0 5731 122
rect 5989 0 6045 122
rect 6287 0 6496 122
rect 6660 0 14387 122
rect 14703 0 14983 122
<< metal3 >>
rect 14438 9997 14785 12893
rect 1680 0 1784 66
rect 3449 0 3782 113
rect 4015 0 4245 282
rect 5787 0 5933 66
rect 14438 0 14652 66
<< obsm3 >>
rect 193 12973 14940 40000
rect 193 9917 14358 12973
rect 14865 9917 14940 12973
rect 193 362 14940 9917
rect 193 193 3935 362
rect 193 146 3369 193
rect 193 66 1600 146
rect 1864 66 3369 146
rect 3862 66 3935 193
rect 4325 146 14940 362
rect 4325 66 5707 146
rect 6013 66 14358 146
rect 14732 66 14940 146
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< obsm4 >>
rect 334 35077 14666 40000
rect 193 19080 14807 35077
rect 334 13927 14666 19080
rect 193 13787 14807 13927
rect 334 12737 14666 13787
rect 193 12617 14807 12737
rect 334 11567 14666 12617
rect 193 11427 14807 11567
rect 334 10349 14666 10545
rect 193 9327 14807 9467
rect 334 8237 14666 9327
rect 193 8117 14807 8237
rect 334 7267 14666 8117
rect 193 7147 14807 7267
rect 334 6297 14666 7147
rect 193 6177 14807 6297
rect 334 5087 14666 6177
rect 193 4967 14807 5087
rect 334 3877 14666 4967
rect 193 3757 14807 3877
rect 273 2907 14727 3757
rect 193 2787 14807 2907
rect 334 1697 14666 2787
rect 193 1577 14807 1697
rect 334 407 14666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 3450 21691 10887 32857
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 7368 15000 8017
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 574 34837 14426 40000
rect 0 33177 15000 34837
rect 0 21371 3130 33177
rect 11207 21371 15000 33177
rect 0 19317 15000 21371
rect 574 3657 14426 19317
rect 513 3007 14487 3657
rect 574 427 14426 3007
<< labels >>
rlabel metal3 s 3449 0 3782 113 6 PAD_A_ESD_H
port 1 nsew signal bidirectional
rlabel metal2 s 3449 0 3782 113 6 PAD_A_ESD_H
port 2 nsew signal bidirectional
rlabel metal3 s 5787 0 5933 66 6 XRES_H_N
port 3 nsew signal output
rlabel metal2 s 5787 0 5933 66 6 XRES_H_N
port 4 nsew signal output
rlabel metal3 s 4015 0 4245 282 6 FILT_IN_H
port 5 nsew signal input
rlabel metal2 s 4015 0 4245 282 6 FILT_IN_H
port 6 nsew signal input
rlabel metal3 s 1680 0 1784 66 6 ENABLE_VDDIO
port 7 nsew signal input
rlabel metal2 s 1685 0 1779 66 6 ENABLE_VDDIO
port 8 nsew signal input
rlabel metal3 s 14438 0 14652 66 6 TIE_WEAK_HI_H
port 9 nsew signal bidirectional
rlabel metal2 s 14443 0 14647 66 6 TIE_WEAK_HI_H
port 10 nsew signal bidirectional
rlabel metal3 s 14438 9997 14785 12893 6 TIE_WEAK_HI_H
port 10 nsew signal bidirectional
rlabel metal2 s 2457 0 2509 66 6 ENABLE_H
port 11 nsew signal input
rlabel metal1 s 2457 0 2509 66 6 ENABLE_H
port 12 nsew signal input
rlabel metal2 s 2911 0 3027 66 6 PULLUP_H
port 13 nsew signal bidirectional
rlabel metal1 s 2911 0 3027 66 6 PULLUP_H
port 14 nsew signal bidirectional
rlabel metal2 s 4472 0 4532 66 6 EN_VDDIO_SIG_H
port 15 nsew signal input
rlabel metal1 s 4472 0 4532 66 6 EN_VDDIO_SIG_H
port 16 nsew signal input
rlabel metal2 s 5864 1072 5916 2217 6 EN_VDDIO_SIG_H
port 16 nsew signal input
rlabel metal2 s 5516 0 5646 66 6 TIE_LO_ESD
port 17 nsew signal output
rlabel metal1 s 5516 0 5646 66 6 TIE_LO_ESD
port 18 nsew signal output
rlabel metal2 s 6101 0 6231 66 6 TIE_HI_ESD
port 19 nsew signal output
rlabel metal1 s 6101 0 6231 66 6 TIE_HI_ESD
port 20 nsew signal output
rlabel metal2 s 6552 0 6604 66 6 DISABLE_PULLUP_H
port 21 nsew signal input
rlabel metal1 s 6552 0 6604 66 6 DISABLE_PULLUP_H
port 22 nsew signal input
rlabel metal1 s 4981 0 5027 1995 6 INP_SEL_H
port 23 nsew signal input
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 24 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 25 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 26 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 27 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 28 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 29 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 30 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 31 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 31 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 31 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 31 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 31 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 31 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 31 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 32 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 33 nsew ground bidirectional
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 34 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 35 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 36 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 6 VSSA
port 37 nsew ground bidirectional
rlabel metal4 s 0 9547 254 9613 6 VSSA
port 38 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 39 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 41 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 42 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 43 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 43 nsew ground bidirectional
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 43 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 43 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 43 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 43 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 43 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 43 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 43 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 44 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 45 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 46 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 47 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 47 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 47 nsew ground bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 48 nsew signal bidirectional
rlabel metal4 s 0 9673 254 10269 6 AMUXBUS_B
port 49 nsew signal bidirectional
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 50 nsew signal bidirectional
rlabel metal4 s 0 10625 254 11221 6 AMUXBUS_A
port 51 nsew signal bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 52 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 53 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 54 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 55 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 55 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 55 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 56 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 57 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 58 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 59 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 60 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 61 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 62 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 63 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 63 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 63 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 63 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 63 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 63 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 63 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 64 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 65 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 66 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 67 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 67 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 67 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 68 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 69 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 70 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 71 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 71 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 71 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 72 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 73 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 74 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 75 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 75 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 75 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 76 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 77 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 78 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 79 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 79 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 79 nsew power bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 80 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 81 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 82 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 83 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 83 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 83 nsew ground bidirectional
rlabel metal5 s 3450 21691 10887 32857 6 PAD
port 84 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass PAD
string LEFsymmetry R90
string LEFview TRUE
string GDS_END 8022630
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3929258
<< end >>
