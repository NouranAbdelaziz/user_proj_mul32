magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< pwell >>
rect 112 1064 768 1086
rect 0 454 880 1064
rect 112 432 768 454
<< nmos >>
rect 194 458 224 1060
rect 348 458 378 1060
rect 502 458 532 1060
rect 656 458 686 1060
<< ndiff >>
rect 138 1048 194 1060
rect 138 1014 149 1048
rect 183 1014 194 1048
rect 138 980 194 1014
rect 138 946 149 980
rect 183 946 194 980
rect 138 912 194 946
rect 138 878 149 912
rect 183 878 194 912
rect 138 844 194 878
rect 138 810 149 844
rect 183 810 194 844
rect 138 776 194 810
rect 138 742 149 776
rect 183 742 194 776
rect 138 708 194 742
rect 138 674 149 708
rect 183 674 194 708
rect 138 640 194 674
rect 138 606 149 640
rect 183 606 194 640
rect 138 572 194 606
rect 138 538 149 572
rect 183 538 194 572
rect 138 504 194 538
rect 138 470 149 504
rect 183 470 194 504
rect 138 458 194 470
rect 224 1048 348 1060
rect 224 470 235 1048
rect 337 470 348 1048
rect 224 458 348 470
rect 378 1048 502 1060
rect 378 470 389 1048
rect 491 470 502 1048
rect 378 458 502 470
rect 532 1048 656 1060
rect 532 470 543 1048
rect 645 470 656 1048
rect 532 458 656 470
rect 686 1048 742 1060
rect 686 1014 697 1048
rect 731 1014 742 1048
rect 686 980 742 1014
rect 686 946 697 980
rect 731 946 742 980
rect 686 912 742 946
rect 686 878 697 912
rect 731 878 742 912
rect 686 844 742 878
rect 686 810 697 844
rect 731 810 742 844
rect 686 776 742 810
rect 686 742 697 776
rect 731 742 742 776
rect 686 708 742 742
rect 686 674 697 708
rect 731 674 742 708
rect 686 640 742 674
rect 686 606 697 640
rect 731 606 742 640
rect 686 572 742 606
rect 686 538 697 572
rect 731 538 742 572
rect 686 504 742 538
rect 686 470 697 504
rect 731 470 742 504
rect 686 458 742 470
<< ndiffc >>
rect 149 1014 183 1048
rect 149 946 183 980
rect 149 878 183 912
rect 149 810 183 844
rect 149 742 183 776
rect 149 674 183 708
rect 149 606 183 640
rect 149 538 183 572
rect 149 470 183 504
rect 235 470 337 1048
rect 389 470 491 1048
rect 543 470 645 1048
rect 697 1014 731 1048
rect 697 946 731 980
rect 697 878 731 912
rect 697 810 731 844
rect 697 742 731 776
rect 697 674 731 708
rect 697 606 731 640
rect 697 538 731 572
rect 697 470 731 504
<< psubdiff >>
rect 26 1014 84 1038
rect 26 980 38 1014
rect 72 980 84 1014
rect 26 946 84 980
rect 26 912 38 946
rect 72 912 84 946
rect 26 878 84 912
rect 26 844 38 878
rect 72 844 84 878
rect 26 810 84 844
rect 26 776 38 810
rect 72 776 84 810
rect 26 742 84 776
rect 26 708 38 742
rect 72 708 84 742
rect 26 674 84 708
rect 26 640 38 674
rect 72 640 84 674
rect 26 606 84 640
rect 26 572 38 606
rect 72 572 84 606
rect 26 538 84 572
rect 26 504 38 538
rect 72 504 84 538
rect 26 480 84 504
rect 796 1014 854 1038
rect 796 980 808 1014
rect 842 980 854 1014
rect 796 946 854 980
rect 796 912 808 946
rect 842 912 854 946
rect 796 878 854 912
rect 796 844 808 878
rect 842 844 854 878
rect 796 810 854 844
rect 796 776 808 810
rect 842 776 854 810
rect 796 742 854 776
rect 796 708 808 742
rect 842 708 854 742
rect 796 674 854 708
rect 796 640 808 674
rect 842 640 854 674
rect 796 606 854 640
rect 796 572 808 606
rect 842 572 854 606
rect 796 538 854 572
rect 796 504 808 538
rect 842 504 854 538
rect 796 480 854 504
<< psubdiffcont >>
rect 38 980 72 1014
rect 38 912 72 946
rect 38 844 72 878
rect 38 776 72 810
rect 38 708 72 742
rect 38 640 72 674
rect 38 572 72 606
rect 38 504 72 538
rect 808 980 842 1014
rect 808 912 842 946
rect 808 844 842 878
rect 808 776 842 810
rect 808 708 842 742
rect 808 640 842 674
rect 808 572 842 606
rect 808 504 842 538
<< poly >>
rect 168 1142 710 1158
rect 168 1108 184 1142
rect 218 1108 252 1142
rect 286 1108 320 1142
rect 354 1108 388 1142
rect 422 1108 456 1142
rect 490 1108 524 1142
rect 558 1108 592 1142
rect 626 1108 660 1142
rect 694 1108 710 1142
rect 168 1092 710 1108
rect 194 1060 224 1092
rect 348 1060 378 1092
rect 502 1060 532 1092
rect 656 1060 686 1092
rect 194 426 224 458
rect 348 426 378 458
rect 502 426 532 458
rect 656 426 686 458
rect 168 410 710 426
rect 168 376 184 410
rect 218 376 252 410
rect 286 376 320 410
rect 354 376 388 410
rect 422 376 456 410
rect 490 376 524 410
rect 558 376 592 410
rect 626 376 660 410
rect 694 376 710 410
rect 168 360 710 376
<< polycont >>
rect 184 1108 218 1142
rect 252 1108 286 1142
rect 320 1108 354 1142
rect 388 1108 422 1142
rect 456 1108 490 1142
rect 524 1108 558 1142
rect 592 1108 626 1142
rect 660 1108 694 1142
rect 184 376 218 410
rect 252 376 286 410
rect 320 376 354 410
rect 388 376 422 410
rect 456 376 490 410
rect 524 376 558 410
rect 592 376 626 410
rect 660 376 694 410
<< locali >>
rect 22 1014 88 1119
rect 168 1108 170 1142
rect 218 1108 252 1142
rect 300 1108 320 1142
rect 354 1108 362 1142
rect 422 1108 456 1142
rect 492 1108 524 1142
rect 588 1108 592 1142
rect 626 1108 650 1142
rect 694 1108 710 1142
rect 22 958 38 1014
rect 72 958 88 1014
rect 22 946 88 958
rect 22 886 38 946
rect 72 886 88 946
rect 22 878 88 886
rect 22 814 38 878
rect 72 814 88 878
rect 22 810 88 814
rect 22 708 38 810
rect 72 708 88 810
rect 22 704 88 708
rect 22 640 38 704
rect 72 640 88 704
rect 22 632 88 640
rect 22 572 38 632
rect 72 572 88 632
rect 22 560 88 572
rect 22 504 38 560
rect 72 504 88 560
rect 22 399 88 504
rect 138 1048 183 1064
rect 138 1033 149 1048
rect 138 999 147 1033
rect 181 999 183 1014
rect 138 980 183 999
rect 138 961 149 980
rect 138 927 147 961
rect 181 927 183 946
rect 138 912 183 927
rect 138 889 149 912
rect 138 855 147 889
rect 181 855 183 878
rect 138 844 183 855
rect 138 817 149 844
rect 138 783 147 817
rect 181 783 183 810
rect 138 776 183 783
rect 138 745 149 776
rect 138 711 147 745
rect 181 711 183 742
rect 138 708 183 711
rect 138 674 149 708
rect 138 673 183 674
rect 138 639 147 673
rect 181 640 183 673
rect 138 606 149 639
rect 138 601 183 606
rect 138 567 147 601
rect 181 572 183 601
rect 138 538 149 567
rect 138 529 183 538
rect 138 495 147 529
rect 181 504 183 529
rect 138 470 149 495
rect 138 454 183 470
rect 233 1048 339 1064
rect 233 1033 235 1048
rect 337 1033 339 1048
rect 233 470 235 495
rect 337 470 339 495
rect 233 454 339 470
rect 387 1048 493 1064
rect 387 1023 389 1048
rect 491 1023 493 1048
rect 387 470 389 485
rect 491 470 493 485
rect 387 454 493 470
rect 541 1048 647 1064
rect 541 1033 543 1048
rect 645 1033 647 1048
rect 541 470 543 495
rect 645 470 647 495
rect 541 454 647 470
rect 697 1048 742 1064
rect 731 1033 742 1048
rect 697 999 699 1014
rect 733 999 742 1033
rect 697 980 742 999
rect 731 961 742 980
rect 697 927 699 946
rect 733 927 742 961
rect 697 912 742 927
rect 731 889 742 912
rect 697 855 699 878
rect 733 855 742 889
rect 697 844 742 855
rect 731 817 742 844
rect 697 783 699 810
rect 733 783 742 817
rect 697 776 742 783
rect 731 745 742 776
rect 697 711 699 742
rect 733 711 742 745
rect 697 708 742 711
rect 731 674 742 708
rect 697 673 742 674
rect 697 640 699 673
rect 733 639 742 673
rect 731 606 742 639
rect 697 601 742 606
rect 697 572 699 601
rect 733 567 742 601
rect 731 538 742 567
rect 697 529 742 538
rect 697 504 699 529
rect 733 495 742 529
rect 731 470 742 495
rect 697 454 742 470
rect 792 1014 858 1119
rect 792 958 808 1014
rect 842 958 858 1014
rect 792 946 858 958
rect 792 886 808 946
rect 842 886 858 946
rect 792 878 858 886
rect 792 814 808 878
rect 842 814 858 878
rect 792 810 858 814
rect 792 708 808 810
rect 842 708 858 810
rect 792 704 858 708
rect 792 640 808 704
rect 842 640 858 704
rect 792 632 858 640
rect 792 572 808 632
rect 842 572 858 632
rect 792 560 858 572
rect 792 504 808 560
rect 842 504 858 560
rect 168 376 170 410
rect 218 376 252 410
rect 300 376 320 410
rect 354 376 362 410
rect 422 376 456 410
rect 492 376 524 410
rect 588 376 592 410
rect 626 376 650 410
rect 694 376 710 410
rect 792 399 858 504
<< viali >>
rect 170 1108 184 1142
rect 184 1108 204 1142
rect 266 1108 286 1142
rect 286 1108 300 1142
rect 362 1108 388 1142
rect 388 1108 396 1142
rect 458 1108 490 1142
rect 490 1108 492 1142
rect 554 1108 558 1142
rect 558 1108 588 1142
rect 650 1108 660 1142
rect 660 1108 684 1142
rect 38 980 72 992
rect 38 958 72 980
rect 38 912 72 920
rect 38 886 72 912
rect 38 844 72 848
rect 38 814 72 844
rect 38 742 72 776
rect 38 674 72 704
rect 38 670 72 674
rect 38 606 72 632
rect 38 598 72 606
rect 38 538 72 560
rect 38 526 72 538
rect 147 1014 149 1033
rect 149 1014 181 1033
rect 147 999 181 1014
rect 147 946 149 961
rect 149 946 181 961
rect 147 927 181 946
rect 147 878 149 889
rect 149 878 181 889
rect 147 855 181 878
rect 147 810 149 817
rect 149 810 181 817
rect 147 783 181 810
rect 147 742 149 745
rect 149 742 181 745
rect 147 711 181 742
rect 147 640 181 673
rect 147 639 149 640
rect 149 639 181 640
rect 147 572 181 601
rect 147 567 149 572
rect 149 567 181 572
rect 147 504 181 529
rect 147 495 149 504
rect 149 495 181 504
rect 233 495 235 1033
rect 235 495 337 1033
rect 337 495 339 1033
rect 387 485 389 1023
rect 389 485 491 1023
rect 491 485 493 1023
rect 541 495 543 1033
rect 543 495 645 1033
rect 645 495 647 1033
rect 699 1014 731 1033
rect 731 1014 733 1033
rect 699 999 733 1014
rect 699 946 731 961
rect 731 946 733 961
rect 699 927 733 946
rect 699 878 731 889
rect 731 878 733 889
rect 699 855 733 878
rect 699 810 731 817
rect 731 810 733 817
rect 699 783 733 810
rect 699 742 731 745
rect 731 742 733 745
rect 699 711 733 742
rect 699 640 733 673
rect 699 639 731 640
rect 731 639 733 640
rect 699 572 733 601
rect 699 567 731 572
rect 731 567 733 572
rect 699 504 733 529
rect 699 495 731 504
rect 731 495 733 504
rect 808 980 842 992
rect 808 958 842 980
rect 808 912 842 920
rect 808 886 842 912
rect 808 844 842 848
rect 808 814 842 844
rect 808 742 842 776
rect 808 674 842 704
rect 808 670 842 674
rect 808 606 842 632
rect 808 598 842 606
rect 808 538 842 560
rect 808 526 842 538
rect 170 376 184 410
rect 184 376 204 410
rect 266 376 286 410
rect 286 376 300 410
rect 362 376 388 410
rect 388 376 396 410
rect 458 376 490 410
rect 490 376 492 410
rect 554 376 558 410
rect 558 376 588 410
rect 650 376 660 410
rect 660 376 684 410
<< metal1 >>
rect 164 1142 690 1154
rect 164 1108 170 1142
rect 204 1108 266 1142
rect 300 1108 362 1142
rect 396 1108 458 1142
rect 492 1108 554 1142
rect 588 1108 650 1142
rect 684 1108 690 1142
rect 164 1096 690 1108
rect 138 1033 194 1060
rect 138 999 147 1033
rect 181 999 194 1033
rect 26 992 84 998
rect 26 958 38 992
rect 72 958 84 992
rect 26 920 84 958
rect 26 886 38 920
rect 72 886 84 920
rect 26 848 84 886
rect 26 814 38 848
rect 72 814 84 848
rect 26 776 84 814
rect 26 742 38 776
rect 72 742 84 776
rect 26 704 84 742
rect 26 670 38 704
rect 72 670 84 704
rect 26 632 84 670
rect 26 598 38 632
rect 72 598 84 632
rect 26 560 84 598
rect 26 526 38 560
rect 72 526 84 560
rect 26 520 84 526
rect 138 964 194 999
rect 138 912 142 964
rect 138 900 194 912
rect 138 848 142 900
rect 138 836 194 848
rect 138 784 142 836
rect 138 783 147 784
rect 181 783 194 784
rect 138 772 194 783
rect 138 720 142 772
rect 138 711 147 720
rect 181 711 194 720
rect 138 708 194 711
rect 138 656 142 708
rect 138 644 147 656
rect 181 644 194 656
rect 138 592 142 644
rect 138 580 147 592
rect 181 580 194 592
rect 138 528 142 580
rect 138 516 147 528
rect 181 516 194 528
rect 138 464 142 516
rect 138 458 194 464
rect 223 1054 349 1060
rect 223 554 228 1054
rect 344 554 349 1054
rect 223 495 233 554
rect 339 495 349 554
rect 223 458 349 495
rect 377 1023 503 1060
rect 377 964 387 1023
rect 493 964 503 1023
rect 377 464 382 964
rect 498 464 503 964
rect 377 458 503 464
rect 531 1054 657 1060
rect 531 554 536 1054
rect 652 554 657 1054
rect 531 495 541 554
rect 647 495 657 554
rect 531 458 657 495
rect 686 1033 742 1060
rect 686 999 699 1033
rect 733 999 742 1033
rect 686 964 742 999
rect 738 912 742 964
rect 686 900 742 912
rect 738 848 742 900
rect 686 836 742 848
rect 738 784 742 836
rect 686 783 699 784
rect 733 783 742 784
rect 686 772 742 783
rect 738 720 742 772
rect 686 711 699 720
rect 733 711 742 720
rect 686 708 742 711
rect 738 656 742 708
rect 686 644 699 656
rect 733 644 742 656
rect 738 592 742 644
rect 686 580 699 592
rect 733 580 742 592
rect 738 528 742 580
rect 686 516 699 528
rect 733 516 742 528
rect 796 992 854 998
rect 796 958 808 992
rect 842 958 854 992
rect 796 920 854 958
rect 796 886 808 920
rect 842 886 854 920
rect 796 848 854 886
rect 796 814 808 848
rect 842 814 854 848
rect 796 776 854 814
rect 796 742 808 776
rect 842 742 854 776
rect 796 704 854 742
rect 796 670 808 704
rect 842 670 854 704
rect 796 632 854 670
rect 796 598 808 632
rect 842 598 854 632
rect 796 560 854 598
rect 796 526 808 560
rect 842 526 854 560
rect 796 520 854 526
rect 738 464 742 516
rect 686 458 742 464
rect 164 410 690 422
rect 164 376 170 410
rect 204 376 266 410
rect 300 376 362 410
rect 396 376 458 410
rect 492 376 554 410
rect 588 376 650 410
rect 684 376 690 410
rect 164 364 690 376
<< via1 >>
rect 142 961 194 964
rect 142 927 147 961
rect 147 927 181 961
rect 181 927 194 961
rect 142 912 194 927
rect 142 889 194 900
rect 142 855 147 889
rect 147 855 181 889
rect 181 855 194 889
rect 142 848 194 855
rect 142 817 194 836
rect 142 784 147 817
rect 147 784 181 817
rect 181 784 194 817
rect 142 745 194 772
rect 142 720 147 745
rect 147 720 181 745
rect 181 720 194 745
rect 142 673 194 708
rect 142 656 147 673
rect 147 656 181 673
rect 181 656 194 673
rect 142 639 147 644
rect 147 639 181 644
rect 181 639 194 644
rect 142 601 194 639
rect 142 592 147 601
rect 147 592 181 601
rect 181 592 194 601
rect 142 567 147 580
rect 147 567 181 580
rect 181 567 194 580
rect 142 529 194 567
rect 142 528 147 529
rect 147 528 181 529
rect 181 528 194 529
rect 142 495 147 516
rect 147 495 181 516
rect 181 495 194 516
rect 142 464 194 495
rect 228 1033 344 1054
rect 228 554 233 1033
rect 233 554 339 1033
rect 339 554 344 1033
rect 382 485 387 964
rect 387 485 493 964
rect 493 485 498 964
rect 382 464 498 485
rect 536 1033 652 1054
rect 536 554 541 1033
rect 541 554 647 1033
rect 647 554 652 1033
rect 686 961 738 964
rect 686 927 699 961
rect 699 927 733 961
rect 733 927 738 961
rect 686 912 738 927
rect 686 889 738 900
rect 686 855 699 889
rect 699 855 733 889
rect 733 855 738 889
rect 686 848 738 855
rect 686 817 738 836
rect 686 784 699 817
rect 699 784 733 817
rect 733 784 738 817
rect 686 745 738 772
rect 686 720 699 745
rect 699 720 733 745
rect 733 720 738 745
rect 686 673 738 708
rect 686 656 699 673
rect 699 656 733 673
rect 733 656 738 673
rect 686 639 699 644
rect 699 639 733 644
rect 733 639 738 644
rect 686 601 738 639
rect 686 592 699 601
rect 699 592 733 601
rect 733 592 738 601
rect 686 567 699 580
rect 699 567 733 580
rect 733 567 738 580
rect 686 529 738 567
rect 686 528 699 529
rect 699 528 733 529
rect 733 528 738 529
rect 686 495 699 516
rect 699 495 733 516
rect 733 495 738 516
rect 686 464 738 495
<< metal2 >>
rect 0 1054 880 1518
rect 0 998 228 1054
rect 112 964 194 970
rect 112 912 142 964
rect 112 900 194 912
rect 112 848 142 900
rect 112 836 194 848
rect 112 784 142 836
rect 112 772 194 784
rect 112 720 142 772
rect 112 708 194 720
rect 112 656 142 708
rect 112 644 194 656
rect 112 592 142 644
rect 112 580 194 592
rect 112 528 142 580
rect 223 554 228 998
rect 344 998 536 1054
rect 344 554 349 998
rect 223 548 349 554
rect 377 964 503 970
rect 112 520 194 528
rect 377 520 382 964
rect 0 516 382 520
rect 0 464 142 516
rect 194 464 382 516
rect 498 520 503 964
rect 531 554 536 998
rect 652 998 880 1054
rect 652 554 657 998
rect 531 548 657 554
rect 686 964 768 970
rect 738 912 768 964
rect 686 900 768 912
rect 738 848 768 900
rect 686 836 768 848
rect 738 784 768 836
rect 686 772 768 784
rect 738 720 768 772
rect 686 708 768 720
rect 738 656 768 708
rect 686 644 768 656
rect 738 592 768 644
rect 686 580 768 592
rect 738 528 768 580
rect 686 520 768 528
rect 498 516 880 520
rect 498 464 686 516
rect 738 464 880 516
rect 0 0 880 464
<< labels >>
flabel comment s 584 762 584 762 0 FreeSans 300 0 0 0 D
flabel comment s 714 745 714 745 0 FreeSans 300 180 0 0 S
flabel comment s 436 762 436 762 0 FreeSans 300 0 0 0 S
flabel comment s 276 762 276 762 0 FreeSans 300 0 0 0 D
flabel comment s 166 745 166 745 0 FreeSans 300 0 0 0 S
flabel metal1 s 36 726 62 793 0 FreeSans 400 90 0 0 SUBSTRATE
flabel metal1 s 416 378 502 403 0 FreeSans 400 0 0 0 GATE
flabel metal2 s 88 22 164 47 0 FreeSans 400 0 0 0 SOURCE
flabel metal2 s 84 1471 173 1503 0 FreeSans 400 0 0 0 DRAIN
<< properties >>
string GDS_END 3164804
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3142608
<< end >>
