magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal3 >>
rect 12409 34239 14940 39600
rect 10151 11248 14858 12136
rect 100 4768 4880 5696
rect 10151 4768 14858 5696
<< obsm3 >>
rect 100 11248 4880 39600
<< metal4 >>
rect 0 39594 254 39600
rect 0 34767 2580 39594
rect 0 34757 254 34767
rect 14746 39594 15000 39600
rect 12415 34767 15000 39594
rect 14746 34757 15000 34767
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 270 12070 334 12134
rect 352 12070 416 12134
rect 434 12070 498 12134
rect 516 12070 580 12134
rect 598 12070 662 12134
rect 679 12070 743 12134
rect 760 12070 824 12134
rect 841 12070 905 12134
rect 922 12070 986 12134
rect 1003 12070 1067 12134
rect 1084 12070 1148 12134
rect 1165 12070 1229 12134
rect 1246 12070 1310 12134
rect 1327 12070 1391 12134
rect 1408 12070 1472 12134
rect 1489 12070 1553 12134
rect 1570 12070 1634 12134
rect 1651 12070 1715 12134
rect 1732 12070 1796 12134
rect 1813 12070 1877 12134
rect 1894 12070 1958 12134
rect 1975 12070 2039 12134
rect 2056 12070 2120 12134
rect 2137 12070 2201 12134
rect 2218 12070 2282 12134
rect 2299 12070 2363 12134
rect 2380 12070 2444 12134
rect 2461 12070 2525 12134
rect 2542 12070 2606 12134
rect 2623 12070 2687 12134
rect 2704 12070 2768 12134
rect 2785 12070 2849 12134
rect 2866 12070 2930 12134
rect 2947 12070 3011 12134
rect 3028 12070 3092 12134
rect 3109 12070 3173 12134
rect 3190 12070 3254 12134
rect 3271 12070 3335 12134
rect 3352 12070 3416 12134
rect 3433 12070 3497 12134
rect 3514 12070 3578 12134
rect 3595 12070 3659 12134
rect 3676 12070 3740 12134
rect 3757 12070 3821 12134
rect 3838 12070 3902 12134
rect 3919 12070 3983 12134
rect 4000 12070 4064 12134
rect 4081 12070 4145 12134
rect 4162 12070 4226 12134
rect 4243 12070 4307 12134
rect 4324 12070 4388 12134
rect 4405 12070 4469 12134
rect 4486 12070 4550 12134
rect 4567 12070 4631 12134
rect 4648 12070 4712 12134
rect 4729 12070 4793 12134
rect 4810 12070 4874 12134
rect 270 11988 334 12052
rect 352 11988 416 12052
rect 434 11988 498 12052
rect 516 11988 580 12052
rect 598 11988 662 12052
rect 679 11988 743 12052
rect 760 11988 824 12052
rect 841 11988 905 12052
rect 922 11988 986 12052
rect 1003 11988 1067 12052
rect 1084 11988 1148 12052
rect 1165 11988 1229 12052
rect 1246 11988 1310 12052
rect 1327 11988 1391 12052
rect 1408 11988 1472 12052
rect 1489 11988 1553 12052
rect 1570 11988 1634 12052
rect 1651 11988 1715 12052
rect 1732 11988 1796 12052
rect 1813 11988 1877 12052
rect 1894 11988 1958 12052
rect 1975 11988 2039 12052
rect 2056 11988 2120 12052
rect 2137 11988 2201 12052
rect 2218 11988 2282 12052
rect 2299 11988 2363 12052
rect 2380 11988 2444 12052
rect 2461 11988 2525 12052
rect 2542 11988 2606 12052
rect 2623 11988 2687 12052
rect 2704 11988 2768 12052
rect 2785 11988 2849 12052
rect 2866 11988 2930 12052
rect 2947 11988 3011 12052
rect 3028 11988 3092 12052
rect 3109 11988 3173 12052
rect 3190 11988 3254 12052
rect 3271 11988 3335 12052
rect 3352 11988 3416 12052
rect 3433 11988 3497 12052
rect 3514 11988 3578 12052
rect 3595 11988 3659 12052
rect 3676 11988 3740 12052
rect 3757 11988 3821 12052
rect 3838 11988 3902 12052
rect 3919 11988 3983 12052
rect 4000 11988 4064 12052
rect 4081 11988 4145 12052
rect 4162 11988 4226 12052
rect 4243 11988 4307 12052
rect 4324 11988 4388 12052
rect 4405 11988 4469 12052
rect 4486 11988 4550 12052
rect 4567 11988 4631 12052
rect 4648 11988 4712 12052
rect 4729 11988 4793 12052
rect 4810 11988 4874 12052
rect 270 11906 334 11970
rect 352 11906 416 11970
rect 434 11906 498 11970
rect 516 11906 580 11970
rect 598 11906 662 11970
rect 679 11906 743 11970
rect 760 11906 824 11970
rect 841 11906 905 11970
rect 922 11906 986 11970
rect 1003 11906 1067 11970
rect 1084 11906 1148 11970
rect 1165 11906 1229 11970
rect 1246 11906 1310 11970
rect 1327 11906 1391 11970
rect 1408 11906 1472 11970
rect 1489 11906 1553 11970
rect 1570 11906 1634 11970
rect 1651 11906 1715 11970
rect 1732 11906 1796 11970
rect 1813 11906 1877 11970
rect 1894 11906 1958 11970
rect 1975 11906 2039 11970
rect 2056 11906 2120 11970
rect 2137 11906 2201 11970
rect 2218 11906 2282 11970
rect 2299 11906 2363 11970
rect 2380 11906 2444 11970
rect 2461 11906 2525 11970
rect 2542 11906 2606 11970
rect 2623 11906 2687 11970
rect 2704 11906 2768 11970
rect 2785 11906 2849 11970
rect 2866 11906 2930 11970
rect 2947 11906 3011 11970
rect 3028 11906 3092 11970
rect 3109 11906 3173 11970
rect 3190 11906 3254 11970
rect 3271 11906 3335 11970
rect 3352 11906 3416 11970
rect 3433 11906 3497 11970
rect 3514 11906 3578 11970
rect 3595 11906 3659 11970
rect 3676 11906 3740 11970
rect 3757 11906 3821 11970
rect 3838 11906 3902 11970
rect 3919 11906 3983 11970
rect 4000 11906 4064 11970
rect 4081 11906 4145 11970
rect 4162 11906 4226 11970
rect 4243 11906 4307 11970
rect 4324 11906 4388 11970
rect 4405 11906 4469 11970
rect 4486 11906 4550 11970
rect 4567 11906 4631 11970
rect 4648 11906 4712 11970
rect 4729 11906 4793 11970
rect 4810 11906 4874 11970
rect 270 11824 334 11888
rect 352 11824 416 11888
rect 434 11824 498 11888
rect 516 11824 580 11888
rect 598 11824 662 11888
rect 679 11824 743 11888
rect 760 11824 824 11888
rect 841 11824 905 11888
rect 922 11824 986 11888
rect 1003 11824 1067 11888
rect 1084 11824 1148 11888
rect 1165 11824 1229 11888
rect 1246 11824 1310 11888
rect 1327 11824 1391 11888
rect 1408 11824 1472 11888
rect 1489 11824 1553 11888
rect 1570 11824 1634 11888
rect 1651 11824 1715 11888
rect 1732 11824 1796 11888
rect 1813 11824 1877 11888
rect 1894 11824 1958 11888
rect 1975 11824 2039 11888
rect 2056 11824 2120 11888
rect 2137 11824 2201 11888
rect 2218 11824 2282 11888
rect 2299 11824 2363 11888
rect 2380 11824 2444 11888
rect 2461 11824 2525 11888
rect 2542 11824 2606 11888
rect 2623 11824 2687 11888
rect 2704 11824 2768 11888
rect 2785 11824 2849 11888
rect 2866 11824 2930 11888
rect 2947 11824 3011 11888
rect 3028 11824 3092 11888
rect 3109 11824 3173 11888
rect 3190 11824 3254 11888
rect 3271 11824 3335 11888
rect 3352 11824 3416 11888
rect 3433 11824 3497 11888
rect 3514 11824 3578 11888
rect 3595 11824 3659 11888
rect 3676 11824 3740 11888
rect 3757 11824 3821 11888
rect 3838 11824 3902 11888
rect 3919 11824 3983 11888
rect 4000 11824 4064 11888
rect 4081 11824 4145 11888
rect 4162 11824 4226 11888
rect 4243 11824 4307 11888
rect 4324 11824 4388 11888
rect 4405 11824 4469 11888
rect 4486 11824 4550 11888
rect 4567 11824 4631 11888
rect 4648 11824 4712 11888
rect 4729 11824 4793 11888
rect 4810 11824 4874 11888
rect 270 11742 334 11806
rect 352 11742 416 11806
rect 434 11742 498 11806
rect 516 11742 580 11806
rect 598 11742 662 11806
rect 679 11742 743 11806
rect 760 11742 824 11806
rect 841 11742 905 11806
rect 922 11742 986 11806
rect 1003 11742 1067 11806
rect 1084 11742 1148 11806
rect 1165 11742 1229 11806
rect 1246 11742 1310 11806
rect 1327 11742 1391 11806
rect 1408 11742 1472 11806
rect 1489 11742 1553 11806
rect 1570 11742 1634 11806
rect 1651 11742 1715 11806
rect 1732 11742 1796 11806
rect 1813 11742 1877 11806
rect 1894 11742 1958 11806
rect 1975 11742 2039 11806
rect 2056 11742 2120 11806
rect 2137 11742 2201 11806
rect 2218 11742 2282 11806
rect 2299 11742 2363 11806
rect 2380 11742 2444 11806
rect 2461 11742 2525 11806
rect 2542 11742 2606 11806
rect 2623 11742 2687 11806
rect 2704 11742 2768 11806
rect 2785 11742 2849 11806
rect 2866 11742 2930 11806
rect 2947 11742 3011 11806
rect 3028 11742 3092 11806
rect 3109 11742 3173 11806
rect 3190 11742 3254 11806
rect 3271 11742 3335 11806
rect 3352 11742 3416 11806
rect 3433 11742 3497 11806
rect 3514 11742 3578 11806
rect 3595 11742 3659 11806
rect 3676 11742 3740 11806
rect 3757 11742 3821 11806
rect 3838 11742 3902 11806
rect 3919 11742 3983 11806
rect 4000 11742 4064 11806
rect 4081 11742 4145 11806
rect 4162 11742 4226 11806
rect 4243 11742 4307 11806
rect 4324 11742 4388 11806
rect 4405 11742 4469 11806
rect 4486 11742 4550 11806
rect 4567 11742 4631 11806
rect 4648 11742 4712 11806
rect 4729 11742 4793 11806
rect 4810 11742 4874 11806
rect 270 11660 334 11724
rect 352 11660 416 11724
rect 434 11660 498 11724
rect 516 11660 580 11724
rect 598 11660 662 11724
rect 679 11660 743 11724
rect 760 11660 824 11724
rect 841 11660 905 11724
rect 922 11660 986 11724
rect 1003 11660 1067 11724
rect 1084 11660 1148 11724
rect 1165 11660 1229 11724
rect 1246 11660 1310 11724
rect 1327 11660 1391 11724
rect 1408 11660 1472 11724
rect 1489 11660 1553 11724
rect 1570 11660 1634 11724
rect 1651 11660 1715 11724
rect 1732 11660 1796 11724
rect 1813 11660 1877 11724
rect 1894 11660 1958 11724
rect 1975 11660 2039 11724
rect 2056 11660 2120 11724
rect 2137 11660 2201 11724
rect 2218 11660 2282 11724
rect 2299 11660 2363 11724
rect 2380 11660 2444 11724
rect 2461 11660 2525 11724
rect 2542 11660 2606 11724
rect 2623 11660 2687 11724
rect 2704 11660 2768 11724
rect 2785 11660 2849 11724
rect 2866 11660 2930 11724
rect 2947 11660 3011 11724
rect 3028 11660 3092 11724
rect 3109 11660 3173 11724
rect 3190 11660 3254 11724
rect 3271 11660 3335 11724
rect 3352 11660 3416 11724
rect 3433 11660 3497 11724
rect 3514 11660 3578 11724
rect 3595 11660 3659 11724
rect 3676 11660 3740 11724
rect 3757 11660 3821 11724
rect 3838 11660 3902 11724
rect 3919 11660 3983 11724
rect 4000 11660 4064 11724
rect 4081 11660 4145 11724
rect 4162 11660 4226 11724
rect 4243 11660 4307 11724
rect 4324 11660 4388 11724
rect 4405 11660 4469 11724
rect 4486 11660 4550 11724
rect 4567 11660 4631 11724
rect 4648 11660 4712 11724
rect 4729 11660 4793 11724
rect 4810 11660 4874 11724
rect 270 11578 334 11642
rect 352 11578 416 11642
rect 434 11578 498 11642
rect 516 11578 580 11642
rect 598 11578 662 11642
rect 679 11578 743 11642
rect 760 11578 824 11642
rect 841 11578 905 11642
rect 922 11578 986 11642
rect 1003 11578 1067 11642
rect 1084 11578 1148 11642
rect 1165 11578 1229 11642
rect 1246 11578 1310 11642
rect 1327 11578 1391 11642
rect 1408 11578 1472 11642
rect 1489 11578 1553 11642
rect 1570 11578 1634 11642
rect 1651 11578 1715 11642
rect 1732 11578 1796 11642
rect 1813 11578 1877 11642
rect 1894 11578 1958 11642
rect 1975 11578 2039 11642
rect 2056 11578 2120 11642
rect 2137 11578 2201 11642
rect 2218 11578 2282 11642
rect 2299 11578 2363 11642
rect 2380 11578 2444 11642
rect 2461 11578 2525 11642
rect 2542 11578 2606 11642
rect 2623 11578 2687 11642
rect 2704 11578 2768 11642
rect 2785 11578 2849 11642
rect 2866 11578 2930 11642
rect 2947 11578 3011 11642
rect 3028 11578 3092 11642
rect 3109 11578 3173 11642
rect 3190 11578 3254 11642
rect 3271 11578 3335 11642
rect 3352 11578 3416 11642
rect 3433 11578 3497 11642
rect 3514 11578 3578 11642
rect 3595 11578 3659 11642
rect 3676 11578 3740 11642
rect 3757 11578 3821 11642
rect 3838 11578 3902 11642
rect 3919 11578 3983 11642
rect 4000 11578 4064 11642
rect 4081 11578 4145 11642
rect 4162 11578 4226 11642
rect 4243 11578 4307 11642
rect 4324 11578 4388 11642
rect 4405 11578 4469 11642
rect 4486 11578 4550 11642
rect 4567 11578 4631 11642
rect 4648 11578 4712 11642
rect 4729 11578 4793 11642
rect 4810 11578 4874 11642
rect 270 11496 334 11560
rect 352 11496 416 11560
rect 434 11496 498 11560
rect 516 11496 580 11560
rect 598 11496 662 11560
rect 679 11496 743 11560
rect 760 11496 824 11560
rect 841 11496 905 11560
rect 922 11496 986 11560
rect 1003 11496 1067 11560
rect 1084 11496 1148 11560
rect 1165 11496 1229 11560
rect 1246 11496 1310 11560
rect 1327 11496 1391 11560
rect 1408 11496 1472 11560
rect 1489 11496 1553 11560
rect 1570 11496 1634 11560
rect 1651 11496 1715 11560
rect 1732 11496 1796 11560
rect 1813 11496 1877 11560
rect 1894 11496 1958 11560
rect 1975 11496 2039 11560
rect 2056 11496 2120 11560
rect 2137 11496 2201 11560
rect 2218 11496 2282 11560
rect 2299 11496 2363 11560
rect 2380 11496 2444 11560
rect 2461 11496 2525 11560
rect 2542 11496 2606 11560
rect 2623 11496 2687 11560
rect 2704 11496 2768 11560
rect 2785 11496 2849 11560
rect 2866 11496 2930 11560
rect 2947 11496 3011 11560
rect 3028 11496 3092 11560
rect 3109 11496 3173 11560
rect 3190 11496 3254 11560
rect 3271 11496 3335 11560
rect 3352 11496 3416 11560
rect 3433 11496 3497 11560
rect 3514 11496 3578 11560
rect 3595 11496 3659 11560
rect 3676 11496 3740 11560
rect 3757 11496 3821 11560
rect 3838 11496 3902 11560
rect 3919 11496 3983 11560
rect 4000 11496 4064 11560
rect 4081 11496 4145 11560
rect 4162 11496 4226 11560
rect 4243 11496 4307 11560
rect 4324 11496 4388 11560
rect 4405 11496 4469 11560
rect 4486 11496 4550 11560
rect 4567 11496 4631 11560
rect 4648 11496 4712 11560
rect 4729 11496 4793 11560
rect 4810 11496 4874 11560
rect 270 11414 334 11478
rect 352 11414 416 11478
rect 434 11414 498 11478
rect 516 11414 580 11478
rect 598 11414 662 11478
rect 679 11414 743 11478
rect 760 11414 824 11478
rect 841 11414 905 11478
rect 922 11414 986 11478
rect 1003 11414 1067 11478
rect 1084 11414 1148 11478
rect 1165 11414 1229 11478
rect 1246 11414 1310 11478
rect 1327 11414 1391 11478
rect 1408 11414 1472 11478
rect 1489 11414 1553 11478
rect 1570 11414 1634 11478
rect 1651 11414 1715 11478
rect 1732 11414 1796 11478
rect 1813 11414 1877 11478
rect 1894 11414 1958 11478
rect 1975 11414 2039 11478
rect 2056 11414 2120 11478
rect 2137 11414 2201 11478
rect 2218 11414 2282 11478
rect 2299 11414 2363 11478
rect 2380 11414 2444 11478
rect 2461 11414 2525 11478
rect 2542 11414 2606 11478
rect 2623 11414 2687 11478
rect 2704 11414 2768 11478
rect 2785 11414 2849 11478
rect 2866 11414 2930 11478
rect 2947 11414 3011 11478
rect 3028 11414 3092 11478
rect 3109 11414 3173 11478
rect 3190 11414 3254 11478
rect 3271 11414 3335 11478
rect 3352 11414 3416 11478
rect 3433 11414 3497 11478
rect 3514 11414 3578 11478
rect 3595 11414 3659 11478
rect 3676 11414 3740 11478
rect 3757 11414 3821 11478
rect 3838 11414 3902 11478
rect 3919 11414 3983 11478
rect 4000 11414 4064 11478
rect 4081 11414 4145 11478
rect 4162 11414 4226 11478
rect 4243 11414 4307 11478
rect 4324 11414 4388 11478
rect 4405 11414 4469 11478
rect 4486 11414 4550 11478
rect 4567 11414 4631 11478
rect 4648 11414 4712 11478
rect 4729 11414 4793 11478
rect 4810 11414 4874 11478
rect 270 11332 334 11396
rect 352 11332 416 11396
rect 434 11332 498 11396
rect 516 11332 580 11396
rect 598 11332 662 11396
rect 679 11332 743 11396
rect 760 11332 824 11396
rect 841 11332 905 11396
rect 922 11332 986 11396
rect 1003 11332 1067 11396
rect 1084 11332 1148 11396
rect 1165 11332 1229 11396
rect 1246 11332 1310 11396
rect 1327 11332 1391 11396
rect 1408 11332 1472 11396
rect 1489 11332 1553 11396
rect 1570 11332 1634 11396
rect 1651 11332 1715 11396
rect 1732 11332 1796 11396
rect 1813 11332 1877 11396
rect 1894 11332 1958 11396
rect 1975 11332 2039 11396
rect 2056 11332 2120 11396
rect 2137 11332 2201 11396
rect 2218 11332 2282 11396
rect 2299 11332 2363 11396
rect 2380 11332 2444 11396
rect 2461 11332 2525 11396
rect 2542 11332 2606 11396
rect 2623 11332 2687 11396
rect 2704 11332 2768 11396
rect 2785 11332 2849 11396
rect 2866 11332 2930 11396
rect 2947 11332 3011 11396
rect 3028 11332 3092 11396
rect 3109 11332 3173 11396
rect 3190 11332 3254 11396
rect 3271 11332 3335 11396
rect 3352 11332 3416 11396
rect 3433 11332 3497 11396
rect 3514 11332 3578 11396
rect 3595 11332 3659 11396
rect 3676 11332 3740 11396
rect 3757 11332 3821 11396
rect 3838 11332 3902 11396
rect 3919 11332 3983 11396
rect 4000 11332 4064 11396
rect 4081 11332 4145 11396
rect 4162 11332 4226 11396
rect 4243 11332 4307 11396
rect 4324 11332 4388 11396
rect 4405 11332 4469 11396
rect 4486 11332 4550 11396
rect 4567 11332 4631 11396
rect 4648 11332 4712 11396
rect 4729 11332 4793 11396
rect 4810 11332 4874 11396
rect 270 11250 334 11314
rect 352 11250 416 11314
rect 434 11250 498 11314
rect 516 11250 580 11314
rect 598 11250 662 11314
rect 679 11250 743 11314
rect 760 11250 824 11314
rect 841 11250 905 11314
rect 922 11250 986 11314
rect 1003 11250 1067 11314
rect 1084 11250 1148 11314
rect 1165 11250 1229 11314
rect 1246 11250 1310 11314
rect 1327 11250 1391 11314
rect 1408 11250 1472 11314
rect 1489 11250 1553 11314
rect 1570 11250 1634 11314
rect 1651 11250 1715 11314
rect 1732 11250 1796 11314
rect 1813 11250 1877 11314
rect 1894 11250 1958 11314
rect 1975 11250 2039 11314
rect 2056 11250 2120 11314
rect 2137 11250 2201 11314
rect 2218 11250 2282 11314
rect 2299 11250 2363 11314
rect 2380 11250 2444 11314
rect 2461 11250 2525 11314
rect 2542 11250 2606 11314
rect 2623 11250 2687 11314
rect 2704 11250 2768 11314
rect 2785 11250 2849 11314
rect 2866 11250 2930 11314
rect 2947 11250 3011 11314
rect 3028 11250 3092 11314
rect 3109 11250 3173 11314
rect 3190 11250 3254 11314
rect 3271 11250 3335 11314
rect 3352 11250 3416 11314
rect 3433 11250 3497 11314
rect 3514 11250 3578 11314
rect 3595 11250 3659 11314
rect 3676 11250 3740 11314
rect 3757 11250 3821 11314
rect 3838 11250 3902 11314
rect 3919 11250 3983 11314
rect 4000 11250 4064 11314
rect 4081 11250 4145 11314
rect 4162 11250 4226 11314
rect 4243 11250 4307 11314
rect 4324 11250 4388 11314
rect 4405 11250 4469 11314
rect 4486 11250 4550 11314
rect 4567 11250 4631 11314
rect 4648 11250 4712 11314
rect 4729 11250 4793 11314
rect 4810 11250 4874 11314
rect 10156 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 10156 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 2660 34687 12335 39600
rect 334 34677 14666 34687
rect 193 18680 14807 34677
rect 334 13527 14666 18680
rect 193 13387 14807 13527
rect 334 12337 14666 13387
rect 193 12217 14807 12337
rect 334 12134 10076 12217
rect 334 12070 352 12134
rect 416 12070 434 12134
rect 498 12070 516 12134
rect 580 12070 598 12134
rect 662 12070 679 12134
rect 743 12070 760 12134
rect 824 12070 841 12134
rect 905 12070 922 12134
rect 986 12070 1003 12134
rect 1067 12070 1084 12134
rect 1148 12070 1165 12134
rect 1229 12070 1246 12134
rect 1310 12070 1327 12134
rect 1391 12070 1408 12134
rect 1472 12070 1489 12134
rect 1553 12070 1570 12134
rect 1634 12070 1651 12134
rect 1715 12070 1732 12134
rect 1796 12070 1813 12134
rect 1877 12070 1894 12134
rect 1958 12070 1975 12134
rect 2039 12070 2056 12134
rect 2120 12070 2137 12134
rect 2201 12070 2218 12134
rect 2282 12070 2299 12134
rect 2363 12070 2380 12134
rect 2444 12070 2461 12134
rect 2525 12070 2542 12134
rect 2606 12070 2623 12134
rect 2687 12070 2704 12134
rect 2768 12070 2785 12134
rect 2849 12070 2866 12134
rect 2930 12070 2947 12134
rect 3011 12070 3028 12134
rect 3092 12070 3109 12134
rect 3173 12070 3190 12134
rect 3254 12070 3271 12134
rect 3335 12070 3352 12134
rect 3416 12070 3433 12134
rect 3497 12070 3514 12134
rect 3578 12070 3595 12134
rect 3659 12070 3676 12134
rect 3740 12070 3757 12134
rect 3821 12070 3838 12134
rect 3902 12070 3919 12134
rect 3983 12070 4000 12134
rect 4064 12070 4081 12134
rect 4145 12070 4162 12134
rect 4226 12070 4243 12134
rect 4307 12070 4324 12134
rect 4388 12070 4405 12134
rect 4469 12070 4486 12134
rect 4550 12070 4567 12134
rect 4631 12070 4648 12134
rect 4712 12070 4729 12134
rect 4793 12070 4810 12134
rect 4874 12070 10076 12134
rect 334 12052 10076 12070
rect 334 11988 352 12052
rect 416 11988 434 12052
rect 498 11988 516 12052
rect 580 11988 598 12052
rect 662 11988 679 12052
rect 743 11988 760 12052
rect 824 11988 841 12052
rect 905 11988 922 12052
rect 986 11988 1003 12052
rect 1067 11988 1084 12052
rect 1148 11988 1165 12052
rect 1229 11988 1246 12052
rect 1310 11988 1327 12052
rect 1391 11988 1408 12052
rect 1472 11988 1489 12052
rect 1553 11988 1570 12052
rect 1634 11988 1651 12052
rect 1715 11988 1732 12052
rect 1796 11988 1813 12052
rect 1877 11988 1894 12052
rect 1958 11988 1975 12052
rect 2039 11988 2056 12052
rect 2120 11988 2137 12052
rect 2201 11988 2218 12052
rect 2282 11988 2299 12052
rect 2363 11988 2380 12052
rect 2444 11988 2461 12052
rect 2525 11988 2542 12052
rect 2606 11988 2623 12052
rect 2687 11988 2704 12052
rect 2768 11988 2785 12052
rect 2849 11988 2866 12052
rect 2930 11988 2947 12052
rect 3011 11988 3028 12052
rect 3092 11988 3109 12052
rect 3173 11988 3190 12052
rect 3254 11988 3271 12052
rect 3335 11988 3352 12052
rect 3416 11988 3433 12052
rect 3497 11988 3514 12052
rect 3578 11988 3595 12052
rect 3659 11988 3676 12052
rect 3740 11988 3757 12052
rect 3821 11988 3838 12052
rect 3902 11988 3919 12052
rect 3983 11988 4000 12052
rect 4064 11988 4081 12052
rect 4145 11988 4162 12052
rect 4226 11988 4243 12052
rect 4307 11988 4324 12052
rect 4388 11988 4405 12052
rect 4469 11988 4486 12052
rect 4550 11988 4567 12052
rect 4631 11988 4648 12052
rect 4712 11988 4729 12052
rect 4793 11988 4810 12052
rect 4874 11988 10076 12052
rect 334 11970 10076 11988
rect 334 11906 352 11970
rect 416 11906 434 11970
rect 498 11906 516 11970
rect 580 11906 598 11970
rect 662 11906 679 11970
rect 743 11906 760 11970
rect 824 11906 841 11970
rect 905 11906 922 11970
rect 986 11906 1003 11970
rect 1067 11906 1084 11970
rect 1148 11906 1165 11970
rect 1229 11906 1246 11970
rect 1310 11906 1327 11970
rect 1391 11906 1408 11970
rect 1472 11906 1489 11970
rect 1553 11906 1570 11970
rect 1634 11906 1651 11970
rect 1715 11906 1732 11970
rect 1796 11906 1813 11970
rect 1877 11906 1894 11970
rect 1958 11906 1975 11970
rect 2039 11906 2056 11970
rect 2120 11906 2137 11970
rect 2201 11906 2218 11970
rect 2282 11906 2299 11970
rect 2363 11906 2380 11970
rect 2444 11906 2461 11970
rect 2525 11906 2542 11970
rect 2606 11906 2623 11970
rect 2687 11906 2704 11970
rect 2768 11906 2785 11970
rect 2849 11906 2866 11970
rect 2930 11906 2947 11970
rect 3011 11906 3028 11970
rect 3092 11906 3109 11970
rect 3173 11906 3190 11970
rect 3254 11906 3271 11970
rect 3335 11906 3352 11970
rect 3416 11906 3433 11970
rect 3497 11906 3514 11970
rect 3578 11906 3595 11970
rect 3659 11906 3676 11970
rect 3740 11906 3757 11970
rect 3821 11906 3838 11970
rect 3902 11906 3919 11970
rect 3983 11906 4000 11970
rect 4064 11906 4081 11970
rect 4145 11906 4162 11970
rect 4226 11906 4243 11970
rect 4307 11906 4324 11970
rect 4388 11906 4405 11970
rect 4469 11906 4486 11970
rect 4550 11906 4567 11970
rect 4631 11906 4648 11970
rect 4712 11906 4729 11970
rect 4793 11906 4810 11970
rect 4874 11906 10076 11970
rect 334 11888 10076 11906
rect 334 11824 352 11888
rect 416 11824 434 11888
rect 498 11824 516 11888
rect 580 11824 598 11888
rect 662 11824 679 11888
rect 743 11824 760 11888
rect 824 11824 841 11888
rect 905 11824 922 11888
rect 986 11824 1003 11888
rect 1067 11824 1084 11888
rect 1148 11824 1165 11888
rect 1229 11824 1246 11888
rect 1310 11824 1327 11888
rect 1391 11824 1408 11888
rect 1472 11824 1489 11888
rect 1553 11824 1570 11888
rect 1634 11824 1651 11888
rect 1715 11824 1732 11888
rect 1796 11824 1813 11888
rect 1877 11824 1894 11888
rect 1958 11824 1975 11888
rect 2039 11824 2056 11888
rect 2120 11824 2137 11888
rect 2201 11824 2218 11888
rect 2282 11824 2299 11888
rect 2363 11824 2380 11888
rect 2444 11824 2461 11888
rect 2525 11824 2542 11888
rect 2606 11824 2623 11888
rect 2687 11824 2704 11888
rect 2768 11824 2785 11888
rect 2849 11824 2866 11888
rect 2930 11824 2947 11888
rect 3011 11824 3028 11888
rect 3092 11824 3109 11888
rect 3173 11824 3190 11888
rect 3254 11824 3271 11888
rect 3335 11824 3352 11888
rect 3416 11824 3433 11888
rect 3497 11824 3514 11888
rect 3578 11824 3595 11888
rect 3659 11824 3676 11888
rect 3740 11824 3757 11888
rect 3821 11824 3838 11888
rect 3902 11824 3919 11888
rect 3983 11824 4000 11888
rect 4064 11824 4081 11888
rect 4145 11824 4162 11888
rect 4226 11824 4243 11888
rect 4307 11824 4324 11888
rect 4388 11824 4405 11888
rect 4469 11824 4486 11888
rect 4550 11824 4567 11888
rect 4631 11824 4648 11888
rect 4712 11824 4729 11888
rect 4793 11824 4810 11888
rect 4874 11824 10076 11888
rect 334 11806 10076 11824
rect 334 11742 352 11806
rect 416 11742 434 11806
rect 498 11742 516 11806
rect 580 11742 598 11806
rect 662 11742 679 11806
rect 743 11742 760 11806
rect 824 11742 841 11806
rect 905 11742 922 11806
rect 986 11742 1003 11806
rect 1067 11742 1084 11806
rect 1148 11742 1165 11806
rect 1229 11742 1246 11806
rect 1310 11742 1327 11806
rect 1391 11742 1408 11806
rect 1472 11742 1489 11806
rect 1553 11742 1570 11806
rect 1634 11742 1651 11806
rect 1715 11742 1732 11806
rect 1796 11742 1813 11806
rect 1877 11742 1894 11806
rect 1958 11742 1975 11806
rect 2039 11742 2056 11806
rect 2120 11742 2137 11806
rect 2201 11742 2218 11806
rect 2282 11742 2299 11806
rect 2363 11742 2380 11806
rect 2444 11742 2461 11806
rect 2525 11742 2542 11806
rect 2606 11742 2623 11806
rect 2687 11742 2704 11806
rect 2768 11742 2785 11806
rect 2849 11742 2866 11806
rect 2930 11742 2947 11806
rect 3011 11742 3028 11806
rect 3092 11742 3109 11806
rect 3173 11742 3190 11806
rect 3254 11742 3271 11806
rect 3335 11742 3352 11806
rect 3416 11742 3433 11806
rect 3497 11742 3514 11806
rect 3578 11742 3595 11806
rect 3659 11742 3676 11806
rect 3740 11742 3757 11806
rect 3821 11742 3838 11806
rect 3902 11742 3919 11806
rect 3983 11742 4000 11806
rect 4064 11742 4081 11806
rect 4145 11742 4162 11806
rect 4226 11742 4243 11806
rect 4307 11742 4324 11806
rect 4388 11742 4405 11806
rect 4469 11742 4486 11806
rect 4550 11742 4567 11806
rect 4631 11742 4648 11806
rect 4712 11742 4729 11806
rect 4793 11742 4810 11806
rect 4874 11742 10076 11806
rect 334 11724 10076 11742
rect 334 11660 352 11724
rect 416 11660 434 11724
rect 498 11660 516 11724
rect 580 11660 598 11724
rect 662 11660 679 11724
rect 743 11660 760 11724
rect 824 11660 841 11724
rect 905 11660 922 11724
rect 986 11660 1003 11724
rect 1067 11660 1084 11724
rect 1148 11660 1165 11724
rect 1229 11660 1246 11724
rect 1310 11660 1327 11724
rect 1391 11660 1408 11724
rect 1472 11660 1489 11724
rect 1553 11660 1570 11724
rect 1634 11660 1651 11724
rect 1715 11660 1732 11724
rect 1796 11660 1813 11724
rect 1877 11660 1894 11724
rect 1958 11660 1975 11724
rect 2039 11660 2056 11724
rect 2120 11660 2137 11724
rect 2201 11660 2218 11724
rect 2282 11660 2299 11724
rect 2363 11660 2380 11724
rect 2444 11660 2461 11724
rect 2525 11660 2542 11724
rect 2606 11660 2623 11724
rect 2687 11660 2704 11724
rect 2768 11660 2785 11724
rect 2849 11660 2866 11724
rect 2930 11660 2947 11724
rect 3011 11660 3028 11724
rect 3092 11660 3109 11724
rect 3173 11660 3190 11724
rect 3254 11660 3271 11724
rect 3335 11660 3352 11724
rect 3416 11660 3433 11724
rect 3497 11660 3514 11724
rect 3578 11660 3595 11724
rect 3659 11660 3676 11724
rect 3740 11660 3757 11724
rect 3821 11660 3838 11724
rect 3902 11660 3919 11724
rect 3983 11660 4000 11724
rect 4064 11660 4081 11724
rect 4145 11660 4162 11724
rect 4226 11660 4243 11724
rect 4307 11660 4324 11724
rect 4388 11660 4405 11724
rect 4469 11660 4486 11724
rect 4550 11660 4567 11724
rect 4631 11660 4648 11724
rect 4712 11660 4729 11724
rect 4793 11660 4810 11724
rect 4874 11660 10076 11724
rect 334 11642 10076 11660
rect 334 11578 352 11642
rect 416 11578 434 11642
rect 498 11578 516 11642
rect 580 11578 598 11642
rect 662 11578 679 11642
rect 743 11578 760 11642
rect 824 11578 841 11642
rect 905 11578 922 11642
rect 986 11578 1003 11642
rect 1067 11578 1084 11642
rect 1148 11578 1165 11642
rect 1229 11578 1246 11642
rect 1310 11578 1327 11642
rect 1391 11578 1408 11642
rect 1472 11578 1489 11642
rect 1553 11578 1570 11642
rect 1634 11578 1651 11642
rect 1715 11578 1732 11642
rect 1796 11578 1813 11642
rect 1877 11578 1894 11642
rect 1958 11578 1975 11642
rect 2039 11578 2056 11642
rect 2120 11578 2137 11642
rect 2201 11578 2218 11642
rect 2282 11578 2299 11642
rect 2363 11578 2380 11642
rect 2444 11578 2461 11642
rect 2525 11578 2542 11642
rect 2606 11578 2623 11642
rect 2687 11578 2704 11642
rect 2768 11578 2785 11642
rect 2849 11578 2866 11642
rect 2930 11578 2947 11642
rect 3011 11578 3028 11642
rect 3092 11578 3109 11642
rect 3173 11578 3190 11642
rect 3254 11578 3271 11642
rect 3335 11578 3352 11642
rect 3416 11578 3433 11642
rect 3497 11578 3514 11642
rect 3578 11578 3595 11642
rect 3659 11578 3676 11642
rect 3740 11578 3757 11642
rect 3821 11578 3838 11642
rect 3902 11578 3919 11642
rect 3983 11578 4000 11642
rect 4064 11578 4081 11642
rect 4145 11578 4162 11642
rect 4226 11578 4243 11642
rect 4307 11578 4324 11642
rect 4388 11578 4405 11642
rect 4469 11578 4486 11642
rect 4550 11578 4567 11642
rect 4631 11578 4648 11642
rect 4712 11578 4729 11642
rect 4793 11578 4810 11642
rect 4874 11578 10076 11642
rect 334 11560 10076 11578
rect 334 11496 352 11560
rect 416 11496 434 11560
rect 498 11496 516 11560
rect 580 11496 598 11560
rect 662 11496 679 11560
rect 743 11496 760 11560
rect 824 11496 841 11560
rect 905 11496 922 11560
rect 986 11496 1003 11560
rect 1067 11496 1084 11560
rect 1148 11496 1165 11560
rect 1229 11496 1246 11560
rect 1310 11496 1327 11560
rect 1391 11496 1408 11560
rect 1472 11496 1489 11560
rect 1553 11496 1570 11560
rect 1634 11496 1651 11560
rect 1715 11496 1732 11560
rect 1796 11496 1813 11560
rect 1877 11496 1894 11560
rect 1958 11496 1975 11560
rect 2039 11496 2056 11560
rect 2120 11496 2137 11560
rect 2201 11496 2218 11560
rect 2282 11496 2299 11560
rect 2363 11496 2380 11560
rect 2444 11496 2461 11560
rect 2525 11496 2542 11560
rect 2606 11496 2623 11560
rect 2687 11496 2704 11560
rect 2768 11496 2785 11560
rect 2849 11496 2866 11560
rect 2930 11496 2947 11560
rect 3011 11496 3028 11560
rect 3092 11496 3109 11560
rect 3173 11496 3190 11560
rect 3254 11496 3271 11560
rect 3335 11496 3352 11560
rect 3416 11496 3433 11560
rect 3497 11496 3514 11560
rect 3578 11496 3595 11560
rect 3659 11496 3676 11560
rect 3740 11496 3757 11560
rect 3821 11496 3838 11560
rect 3902 11496 3919 11560
rect 3983 11496 4000 11560
rect 4064 11496 4081 11560
rect 4145 11496 4162 11560
rect 4226 11496 4243 11560
rect 4307 11496 4324 11560
rect 4388 11496 4405 11560
rect 4469 11496 4486 11560
rect 4550 11496 4567 11560
rect 4631 11496 4648 11560
rect 4712 11496 4729 11560
rect 4793 11496 4810 11560
rect 4874 11496 10076 11560
rect 334 11478 10076 11496
rect 334 11414 352 11478
rect 416 11414 434 11478
rect 498 11414 516 11478
rect 580 11414 598 11478
rect 662 11414 679 11478
rect 743 11414 760 11478
rect 824 11414 841 11478
rect 905 11414 922 11478
rect 986 11414 1003 11478
rect 1067 11414 1084 11478
rect 1148 11414 1165 11478
rect 1229 11414 1246 11478
rect 1310 11414 1327 11478
rect 1391 11414 1408 11478
rect 1472 11414 1489 11478
rect 1553 11414 1570 11478
rect 1634 11414 1651 11478
rect 1715 11414 1732 11478
rect 1796 11414 1813 11478
rect 1877 11414 1894 11478
rect 1958 11414 1975 11478
rect 2039 11414 2056 11478
rect 2120 11414 2137 11478
rect 2201 11414 2218 11478
rect 2282 11414 2299 11478
rect 2363 11414 2380 11478
rect 2444 11414 2461 11478
rect 2525 11414 2542 11478
rect 2606 11414 2623 11478
rect 2687 11414 2704 11478
rect 2768 11414 2785 11478
rect 2849 11414 2866 11478
rect 2930 11414 2947 11478
rect 3011 11414 3028 11478
rect 3092 11414 3109 11478
rect 3173 11414 3190 11478
rect 3254 11414 3271 11478
rect 3335 11414 3352 11478
rect 3416 11414 3433 11478
rect 3497 11414 3514 11478
rect 3578 11414 3595 11478
rect 3659 11414 3676 11478
rect 3740 11414 3757 11478
rect 3821 11414 3838 11478
rect 3902 11414 3919 11478
rect 3983 11414 4000 11478
rect 4064 11414 4081 11478
rect 4145 11414 4162 11478
rect 4226 11414 4243 11478
rect 4307 11414 4324 11478
rect 4388 11414 4405 11478
rect 4469 11414 4486 11478
rect 4550 11414 4567 11478
rect 4631 11414 4648 11478
rect 4712 11414 4729 11478
rect 4793 11414 4810 11478
rect 4874 11414 10076 11478
rect 334 11396 10076 11414
rect 334 11332 352 11396
rect 416 11332 434 11396
rect 498 11332 516 11396
rect 580 11332 598 11396
rect 662 11332 679 11396
rect 743 11332 760 11396
rect 824 11332 841 11396
rect 905 11332 922 11396
rect 986 11332 1003 11396
rect 1067 11332 1084 11396
rect 1148 11332 1165 11396
rect 1229 11332 1246 11396
rect 1310 11332 1327 11396
rect 1391 11332 1408 11396
rect 1472 11332 1489 11396
rect 1553 11332 1570 11396
rect 1634 11332 1651 11396
rect 1715 11332 1732 11396
rect 1796 11332 1813 11396
rect 1877 11332 1894 11396
rect 1958 11332 1975 11396
rect 2039 11332 2056 11396
rect 2120 11332 2137 11396
rect 2201 11332 2218 11396
rect 2282 11332 2299 11396
rect 2363 11332 2380 11396
rect 2444 11332 2461 11396
rect 2525 11332 2542 11396
rect 2606 11332 2623 11396
rect 2687 11332 2704 11396
rect 2768 11332 2785 11396
rect 2849 11332 2866 11396
rect 2930 11332 2947 11396
rect 3011 11332 3028 11396
rect 3092 11332 3109 11396
rect 3173 11332 3190 11396
rect 3254 11332 3271 11396
rect 3335 11332 3352 11396
rect 3416 11332 3433 11396
rect 3497 11332 3514 11396
rect 3578 11332 3595 11396
rect 3659 11332 3676 11396
rect 3740 11332 3757 11396
rect 3821 11332 3838 11396
rect 3902 11332 3919 11396
rect 3983 11332 4000 11396
rect 4064 11332 4081 11396
rect 4145 11332 4162 11396
rect 4226 11332 4243 11396
rect 4307 11332 4324 11396
rect 4388 11332 4405 11396
rect 4469 11332 4486 11396
rect 4550 11332 4567 11396
rect 4631 11332 4648 11396
rect 4712 11332 4729 11396
rect 4793 11332 4810 11396
rect 4874 11332 10076 11396
rect 334 11314 10076 11332
rect 334 11250 352 11314
rect 416 11250 434 11314
rect 498 11250 516 11314
rect 580 11250 598 11314
rect 662 11250 679 11314
rect 743 11250 760 11314
rect 824 11250 841 11314
rect 905 11250 922 11314
rect 986 11250 1003 11314
rect 1067 11250 1084 11314
rect 1148 11250 1165 11314
rect 1229 11250 1246 11314
rect 1310 11250 1327 11314
rect 1391 11250 1408 11314
rect 1472 11250 1489 11314
rect 1553 11250 1570 11314
rect 1634 11250 1651 11314
rect 1715 11250 1732 11314
rect 1796 11250 1813 11314
rect 1877 11250 1894 11314
rect 1958 11250 1975 11314
rect 2039 11250 2056 11314
rect 2120 11250 2137 11314
rect 2201 11250 2218 11314
rect 2282 11250 2299 11314
rect 2363 11250 2380 11314
rect 2444 11250 2461 11314
rect 2525 11250 2542 11314
rect 2606 11250 2623 11314
rect 2687 11250 2704 11314
rect 2768 11250 2785 11314
rect 2849 11250 2866 11314
rect 2930 11250 2947 11314
rect 3011 11250 3028 11314
rect 3092 11250 3109 11314
rect 3173 11250 3190 11314
rect 3254 11250 3271 11314
rect 3335 11250 3352 11314
rect 3416 11250 3433 11314
rect 3497 11250 3514 11314
rect 3578 11250 3595 11314
rect 3659 11250 3676 11314
rect 3740 11250 3757 11314
rect 3821 11250 3838 11314
rect 3902 11250 3919 11314
rect 3983 11250 4000 11314
rect 4064 11250 4081 11314
rect 4145 11250 4162 11314
rect 4226 11250 4243 11314
rect 4307 11250 4324 11314
rect 4388 11250 4405 11314
rect 4469 11250 4486 11314
rect 4550 11250 4567 11314
rect 4631 11250 4648 11314
rect 4712 11250 4729 11314
rect 4793 11250 4810 11314
rect 4874 11250 10076 11314
rect 334 11167 10076 11250
rect 193 11027 14807 11167
rect 334 9949 14666 10145
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 6867 14666 7717
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 10076 5777
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 18917 15000 34437
rect 574 6968 14426 18917
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 10225 254 10821 6 AMUXBUS_A
port 2 nsew signal bidirectional
rlabel metal4 s 14746 10225 15000 10821 6 AMUXBUS_A
port 2 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 3 nsew signal bidirectional
rlabel metal4 s 0 9273 254 9869 6 AMUXBUS_B
port 4 nsew signal bidirectional
rlabel metal4 s 14746 9273 15000 9869 6 AMUXBUS_B
port 4 nsew signal bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 5 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 6 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 12 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 12 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 12 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 13 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 14 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 15 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 16 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 16 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 16 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 16 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 17 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 18 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 19 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 20 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 21 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 22 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 23 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 24 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 24 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 25 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 26 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 27 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 28 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 28 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 28 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 28 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 29 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 31 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 32 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 33 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 34 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 35 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 36 nsew ground bidirectional
rlabel metal4 s 0 9147 254 9213 6 VSSA
port 37 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 38 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 6 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 0 9147 254 9213 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 14746 9147 15000 9213 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 14746 10881 15000 10947 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 41 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 42 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 43 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 44 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 44 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 44 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 44 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 45 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 46 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 47 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 48 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 49 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 50 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 100 4768 4880 5696 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10151 4768 14858 5696 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12409 34239 14940 39600 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 0 39594 254 39600 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 0 34767 2580 39594 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 0 34757 254 34767 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 10156 4767 15000 5697 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 14746 39594 15000 39600 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 34767 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 12415 34767 15000 39594 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 39541 14928 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 39460 14928 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 39379 14928 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 39298 14928 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 39217 14928 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 39136 14928 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 39055 14928 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38974 14928 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38893 14928 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38812 14928 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38731 14928 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38650 14928 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38569 14928 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38488 14928 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38407 14928 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38326 14928 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38245 14928 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38164 14928 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38083 14928 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 38002 14928 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37921 14928 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37840 14928 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37759 14928 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37678 14928 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37597 14928 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37516 14928 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37435 14928 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37354 14928 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37273 14928 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37192 14928 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37111 14928 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 37030 14928 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36949 14928 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36868 14928 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36787 14928 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36706 14928 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36625 14928 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36544 14928 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36463 14928 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36382 14928 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36301 14928 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36220 14928 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36140 14928 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 36060 14928 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35980 14928 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35900 14928 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35820 14928 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35740 14928 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35660 14928 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35580 14928 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35500 14928 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35420 14928 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35340 14928 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35260 14928 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35180 14928 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35100 14928 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 35020 14928 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 34940 14928 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 34860 14928 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14888 34780 14928 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 39541 14846 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 39460 14846 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 39379 14846 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 39298 14846 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 39217 14846 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 39136 14846 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 39055 14846 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38974 14846 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38893 14846 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38812 14846 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38731 14846 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38650 14846 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38569 14846 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38488 14846 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38407 14846 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38326 14846 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38245 14846 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38164 14846 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38083 14846 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 38002 14846 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37921 14846 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37840 14846 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37759 14846 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37678 14846 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37597 14846 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37516 14846 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37435 14846 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37354 14846 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37273 14846 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37192 14846 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37111 14846 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 37030 14846 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36949 14846 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36868 14846 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36787 14846 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36706 14846 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36625 14846 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36544 14846 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36463 14846 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36382 14846 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36301 14846 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36220 14846 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36140 14846 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 36060 14846 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35980 14846 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35900 14846 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35820 14846 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35740 14846 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35660 14846 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35580 14846 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35500 14846 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35420 14846 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35340 14846 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35260 14846 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35180 14846 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35100 14846 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 35020 14846 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 34940 14846 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 34860 14846 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14806 34780 14846 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 5642 14840 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 5556 14840 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 5470 14840 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 5384 14840 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 5298 14840 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 5212 14840 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 5126 14840 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 5040 14840 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 4954 14840 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 4868 14840 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14800 4782 14840 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 39541 14764 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 39460 14764 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 39379 14764 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 39298 14764 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 39217 14764 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 39136 14764 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 39055 14764 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38974 14764 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38893 14764 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38812 14764 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38731 14764 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38650 14764 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38569 14764 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38488 14764 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38407 14764 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38326 14764 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38245 14764 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38164 14764 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38083 14764 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 38002 14764 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37921 14764 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37840 14764 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37759 14764 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37678 14764 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37597 14764 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37516 14764 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37435 14764 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37354 14764 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37273 14764 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37192 14764 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37111 14764 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 37030 14764 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36949 14764 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36868 14764 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36787 14764 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36706 14764 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36625 14764 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36544 14764 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36463 14764 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36382 14764 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36301 14764 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36220 14764 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36140 14764 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 36060 14764 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35980 14764 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35900 14764 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35820 14764 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35740 14764 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35660 14764 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35580 14764 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35500 14764 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35420 14764 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35340 14764 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35260 14764 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35180 14764 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35100 14764 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 35020 14764 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 34940 14764 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 34860 14764 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14724 34780 14764 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 5642 14759 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 5556 14759 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 5470 14759 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 5384 14759 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 5298 14759 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 5212 14759 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 5126 14759 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 5040 14759 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 4954 14759 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 4868 14759 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14719 4782 14759 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 39541 14682 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 39460 14682 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 39379 14682 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 39298 14682 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 39217 14682 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 39136 14682 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 39055 14682 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38974 14682 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38893 14682 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38812 14682 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38731 14682 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38650 14682 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38569 14682 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38488 14682 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38407 14682 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38326 14682 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38245 14682 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38164 14682 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38083 14682 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 38002 14682 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37921 14682 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37840 14682 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37759 14682 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37678 14682 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37597 14682 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37516 14682 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37435 14682 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37354 14682 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37273 14682 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37192 14682 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37111 14682 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 37030 14682 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36949 14682 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36868 14682 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36787 14682 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36706 14682 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36625 14682 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36544 14682 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36463 14682 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36382 14682 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36301 14682 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36220 14682 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36140 14682 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 36060 14682 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35980 14682 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35900 14682 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35820 14682 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35740 14682 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35660 14682 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35580 14682 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35500 14682 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35420 14682 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35340 14682 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35260 14682 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35180 14682 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35100 14682 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 35020 14682 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 34940 14682 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 34860 14682 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14642 34780 14682 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 5642 14678 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 5556 14678 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 5470 14678 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 5384 14678 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 5298 14678 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 5212 14678 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 5126 14678 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 5040 14678 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 4954 14678 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 4868 14678 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14638 4782 14678 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 39541 14600 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 39460 14600 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 39379 14600 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 39298 14600 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 39217 14600 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 39136 14600 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 39055 14600 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38974 14600 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38893 14600 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38812 14600 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38731 14600 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38650 14600 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38569 14600 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38488 14600 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38407 14600 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38326 14600 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38245 14600 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38164 14600 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38083 14600 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 38002 14600 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37921 14600 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37840 14600 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37759 14600 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37678 14600 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37597 14600 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37516 14600 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37435 14600 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37354 14600 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37273 14600 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37192 14600 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37111 14600 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 37030 14600 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36949 14600 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36868 14600 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36787 14600 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36706 14600 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36625 14600 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36544 14600 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36463 14600 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36382 14600 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36301 14600 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36220 14600 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36140 14600 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 36060 14600 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35980 14600 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35900 14600 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35820 14600 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35740 14600 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35660 14600 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35580 14600 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35500 14600 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35420 14600 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35340 14600 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35260 14600 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35180 14600 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35100 14600 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 35020 14600 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 34940 14600 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 34860 14600 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14560 34780 14600 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 5642 14597 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 5556 14597 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 5470 14597 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 5384 14597 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 5298 14597 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 5212 14597 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 5126 14597 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 5040 14597 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 4954 14597 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 4868 14597 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14557 4782 14597 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 39541 14518 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 39460 14518 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 39379 14518 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 39298 14518 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 39217 14518 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 39136 14518 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 39055 14518 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38974 14518 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38893 14518 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38812 14518 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38731 14518 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38650 14518 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38569 14518 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38488 14518 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38407 14518 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38326 14518 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38245 14518 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38164 14518 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38083 14518 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 38002 14518 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37921 14518 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37840 14518 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37759 14518 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37678 14518 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37597 14518 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37516 14518 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37435 14518 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37354 14518 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37273 14518 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37192 14518 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37111 14518 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 37030 14518 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36949 14518 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36868 14518 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36787 14518 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36706 14518 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36625 14518 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36544 14518 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36463 14518 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36382 14518 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36301 14518 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36220 14518 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36140 14518 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 36060 14518 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35980 14518 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35900 14518 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35820 14518 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35740 14518 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35660 14518 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35580 14518 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35500 14518 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35420 14518 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35340 14518 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35260 14518 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35180 14518 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35100 14518 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 35020 14518 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 34940 14518 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 34860 14518 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14478 34780 14518 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 5642 14516 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 5556 14516 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 5470 14516 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 5384 14516 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 5298 14516 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 5212 14516 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 5126 14516 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 5040 14516 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 4954 14516 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 4868 14516 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14476 4782 14516 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 39541 14436 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 39460 14436 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 39379 14436 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 39298 14436 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 39217 14436 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 39136 14436 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 39055 14436 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38974 14436 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38893 14436 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38812 14436 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38731 14436 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38650 14436 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38569 14436 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38488 14436 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38407 14436 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38326 14436 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38245 14436 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38164 14436 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38083 14436 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 38002 14436 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37921 14436 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37840 14436 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37759 14436 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37678 14436 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37597 14436 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37516 14436 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37435 14436 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37354 14436 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37273 14436 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37192 14436 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37111 14436 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 37030 14436 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36949 14436 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36868 14436 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36787 14436 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36706 14436 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36625 14436 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36544 14436 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36463 14436 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36382 14436 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36301 14436 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36220 14436 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36140 14436 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 36060 14436 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35980 14436 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35900 14436 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35820 14436 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35740 14436 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35660 14436 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35580 14436 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35500 14436 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35420 14436 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35340 14436 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35260 14436 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35180 14436 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35100 14436 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 35020 14436 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 34940 14436 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 34860 14436 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14396 34780 14436 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 5642 14435 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 5556 14435 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 5470 14435 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 5384 14435 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 5298 14435 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 5212 14435 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 5126 14435 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 5040 14435 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 4954 14435 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 4868 14435 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14395 4782 14435 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 39541 14354 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 39460 14354 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 39379 14354 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 39298 14354 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 39217 14354 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 39136 14354 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 39055 14354 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38974 14354 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38893 14354 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38812 14354 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38731 14354 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38650 14354 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38569 14354 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38488 14354 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38407 14354 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38326 14354 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38245 14354 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38164 14354 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38083 14354 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 38002 14354 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37921 14354 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37840 14354 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37759 14354 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37678 14354 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37597 14354 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37516 14354 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37435 14354 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37354 14354 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37273 14354 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37192 14354 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37111 14354 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 37030 14354 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36949 14354 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36868 14354 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36787 14354 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36706 14354 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36625 14354 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36544 14354 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36463 14354 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36382 14354 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36301 14354 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36220 14354 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36140 14354 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 36060 14354 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35980 14354 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35900 14354 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35820 14354 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35740 14354 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35660 14354 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35580 14354 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35500 14354 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35420 14354 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35340 14354 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35260 14354 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35180 14354 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35100 14354 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 35020 14354 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 34940 14354 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 34860 14354 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 34780 14354 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 5642 14354 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 5556 14354 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 5470 14354 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 5384 14354 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 5298 14354 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 5212 14354 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 5126 14354 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 5040 14354 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 4954 14354 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 4868 14354 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14314 4782 14354 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 5642 14273 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 5556 14273 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 5470 14273 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 5384 14273 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 5298 14273 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 5212 14273 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 5126 14273 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 5040 14273 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 4954 14273 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 4868 14273 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14233 4782 14273 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 39541 14272 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 39460 14272 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 39379 14272 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 39298 14272 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 39217 14272 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 39136 14272 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 39055 14272 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38974 14272 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38893 14272 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38812 14272 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38731 14272 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38650 14272 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38569 14272 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38488 14272 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38407 14272 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38326 14272 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38245 14272 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38164 14272 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38083 14272 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 38002 14272 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37921 14272 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37840 14272 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37759 14272 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37678 14272 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37597 14272 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37516 14272 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37435 14272 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37354 14272 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37273 14272 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37192 14272 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37111 14272 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 37030 14272 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36949 14272 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36868 14272 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36787 14272 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36706 14272 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36625 14272 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36544 14272 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36463 14272 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36382 14272 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36301 14272 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36220 14272 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36140 14272 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 36060 14272 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35980 14272 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35900 14272 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35820 14272 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35740 14272 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35660 14272 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35580 14272 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35500 14272 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35420 14272 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35340 14272 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35260 14272 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35180 14272 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35100 14272 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 35020 14272 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 34940 14272 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 34860 14272 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14232 34780 14272 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 5642 14192 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 5556 14192 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 5470 14192 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 5384 14192 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 5298 14192 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 5212 14192 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 5126 14192 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 5040 14192 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 4954 14192 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 4868 14192 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14152 4782 14192 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 39541 14190 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 39460 14190 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 39379 14190 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 39298 14190 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 39217 14190 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 39136 14190 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 39055 14190 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38974 14190 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38893 14190 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38812 14190 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38731 14190 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38650 14190 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38569 14190 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38488 14190 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38407 14190 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38326 14190 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38245 14190 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38164 14190 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38083 14190 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 38002 14190 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37921 14190 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37840 14190 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37759 14190 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37678 14190 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37597 14190 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37516 14190 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37435 14190 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37354 14190 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37273 14190 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37192 14190 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37111 14190 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 37030 14190 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36949 14190 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36868 14190 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36787 14190 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36706 14190 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36625 14190 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36544 14190 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36463 14190 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36382 14190 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36301 14190 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36220 14190 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36140 14190 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 36060 14190 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35980 14190 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35900 14190 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35820 14190 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35740 14190 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35660 14190 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35580 14190 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35500 14190 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35420 14190 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35340 14190 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35260 14190 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35180 14190 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35100 14190 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 35020 14190 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 34940 14190 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 34860 14190 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14150 34780 14190 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 5642 14111 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 5556 14111 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 5470 14111 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 5384 14111 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 5298 14111 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 5212 14111 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 5126 14111 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 5040 14111 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 4954 14111 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 4868 14111 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14071 4782 14111 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 39541 14108 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 39460 14108 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 39379 14108 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 39298 14108 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 39217 14108 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 39136 14108 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 39055 14108 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38974 14108 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38893 14108 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38812 14108 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38731 14108 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38650 14108 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38569 14108 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38488 14108 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38407 14108 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38326 14108 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38245 14108 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38164 14108 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38083 14108 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 38002 14108 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37921 14108 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37840 14108 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37759 14108 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37678 14108 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37597 14108 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37516 14108 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37435 14108 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37354 14108 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37273 14108 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37192 14108 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37111 14108 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 37030 14108 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36949 14108 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36868 14108 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36787 14108 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36706 14108 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36625 14108 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36544 14108 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36463 14108 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36382 14108 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36301 14108 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36220 14108 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36140 14108 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 36060 14108 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35980 14108 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35900 14108 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35820 14108 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35740 14108 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35660 14108 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35580 14108 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35500 14108 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35420 14108 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35340 14108 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35260 14108 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35180 14108 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35100 14108 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 35020 14108 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 34940 14108 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 34860 14108 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 14068 34780 14108 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 5642 14030 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 5556 14030 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 5470 14030 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 5384 14030 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 5298 14030 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 5212 14030 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 5126 14030 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 5040 14030 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 4954 14030 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 4868 14030 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13990 4782 14030 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 39541 14026 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 39460 14026 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 39379 14026 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 39298 14026 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 39217 14026 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 39136 14026 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 39055 14026 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38974 14026 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38893 14026 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38812 14026 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38731 14026 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38650 14026 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38569 14026 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38488 14026 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38407 14026 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38326 14026 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38245 14026 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38164 14026 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38083 14026 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 38002 14026 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37921 14026 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37840 14026 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37759 14026 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37678 14026 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37597 14026 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37516 14026 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37435 14026 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37354 14026 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37273 14026 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37192 14026 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37111 14026 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 37030 14026 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36949 14026 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36868 14026 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36787 14026 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36706 14026 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36625 14026 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36544 14026 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36463 14026 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36382 14026 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36301 14026 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36220 14026 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36140 14026 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 36060 14026 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35980 14026 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35900 14026 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35820 14026 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35740 14026 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35660 14026 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35580 14026 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35500 14026 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35420 14026 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35340 14026 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35260 14026 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35180 14026 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35100 14026 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 35020 14026 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 34940 14026 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 34860 14026 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13986 34780 14026 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 5642 13949 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 5556 13949 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 5470 13949 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 5384 13949 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 5298 13949 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 5212 13949 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 5126 13949 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 5040 13949 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 4954 13949 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 4868 13949 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13909 4782 13949 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 39541 13944 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 39460 13944 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 39379 13944 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 39298 13944 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 39217 13944 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 39136 13944 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 39055 13944 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38974 13944 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38893 13944 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38812 13944 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38731 13944 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38650 13944 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38569 13944 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38488 13944 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38407 13944 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38326 13944 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38245 13944 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38164 13944 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38083 13944 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 38002 13944 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37921 13944 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37840 13944 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37759 13944 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37678 13944 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37597 13944 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37516 13944 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37435 13944 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37354 13944 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37273 13944 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37192 13944 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37111 13944 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 37030 13944 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36949 13944 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36868 13944 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36787 13944 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36706 13944 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36625 13944 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36544 13944 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36463 13944 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36382 13944 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36301 13944 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36220 13944 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36140 13944 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 36060 13944 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35980 13944 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35900 13944 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35820 13944 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35740 13944 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35660 13944 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35580 13944 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35500 13944 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35420 13944 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35340 13944 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35260 13944 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35180 13944 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35100 13944 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 35020 13944 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 34940 13944 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 34860 13944 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13904 34780 13944 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 5642 13868 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 5556 13868 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 5470 13868 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 5384 13868 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 5298 13868 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 5212 13868 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 5126 13868 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 5040 13868 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 4954 13868 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 4868 13868 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13828 4782 13868 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 39541 13862 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 39460 13862 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 39379 13862 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 39298 13862 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 39217 13862 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 39136 13862 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 39055 13862 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38974 13862 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38893 13862 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38812 13862 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38731 13862 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38650 13862 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38569 13862 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38488 13862 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38407 13862 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38326 13862 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38245 13862 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38164 13862 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38083 13862 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 38002 13862 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37921 13862 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37840 13862 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37759 13862 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37678 13862 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37597 13862 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37516 13862 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37435 13862 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37354 13862 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37273 13862 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37192 13862 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37111 13862 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 37030 13862 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36949 13862 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36868 13862 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36787 13862 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36706 13862 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36625 13862 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36544 13862 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36463 13862 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36382 13862 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36301 13862 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36220 13862 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36140 13862 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 36060 13862 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35980 13862 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35900 13862 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35820 13862 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35740 13862 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35660 13862 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35580 13862 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35500 13862 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35420 13862 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35340 13862 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35260 13862 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35180 13862 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35100 13862 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 35020 13862 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 34940 13862 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 34860 13862 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13822 34780 13862 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 5642 13787 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 5556 13787 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 5470 13787 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 5384 13787 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 5298 13787 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 5212 13787 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 5126 13787 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 5040 13787 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 4954 13787 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 4868 13787 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13747 4782 13787 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 39541 13780 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 39460 13780 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 39379 13780 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 39298 13780 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 39217 13780 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 39136 13780 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 39055 13780 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38974 13780 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38893 13780 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38812 13780 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38731 13780 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38650 13780 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38569 13780 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38488 13780 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38407 13780 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38326 13780 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38245 13780 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38164 13780 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38083 13780 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 38002 13780 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37921 13780 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37840 13780 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37759 13780 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37678 13780 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37597 13780 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37516 13780 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37435 13780 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37354 13780 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37273 13780 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37192 13780 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37111 13780 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 37030 13780 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36949 13780 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36868 13780 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36787 13780 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36706 13780 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36625 13780 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36544 13780 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36463 13780 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36382 13780 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36301 13780 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36220 13780 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36140 13780 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 36060 13780 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35980 13780 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35900 13780 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35820 13780 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35740 13780 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35660 13780 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35580 13780 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35500 13780 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35420 13780 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35340 13780 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35260 13780 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35180 13780 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35100 13780 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 35020 13780 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 34940 13780 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 34860 13780 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13740 34780 13780 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 5642 13706 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 5556 13706 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 5470 13706 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 5384 13706 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 5298 13706 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 5212 13706 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 5126 13706 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 5040 13706 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 4954 13706 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 4868 13706 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13666 4782 13706 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 39541 13698 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 39460 13698 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 39379 13698 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 39298 13698 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 39217 13698 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 39136 13698 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 39055 13698 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38974 13698 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38893 13698 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38812 13698 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38731 13698 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38650 13698 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38569 13698 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38488 13698 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38407 13698 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38326 13698 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38245 13698 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38164 13698 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38083 13698 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 38002 13698 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37921 13698 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37840 13698 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37759 13698 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37678 13698 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37597 13698 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37516 13698 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37435 13698 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37354 13698 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37273 13698 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37192 13698 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37111 13698 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 37030 13698 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36949 13698 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36868 13698 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36787 13698 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36706 13698 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36625 13698 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36544 13698 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36463 13698 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36382 13698 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36301 13698 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36220 13698 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36140 13698 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 36060 13698 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35980 13698 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35900 13698 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35820 13698 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35740 13698 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35660 13698 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35580 13698 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35500 13698 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35420 13698 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35340 13698 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35260 13698 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35180 13698 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35100 13698 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 35020 13698 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 34940 13698 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 34860 13698 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13658 34780 13698 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 5642 13625 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 5556 13625 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 5470 13625 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 5384 13625 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 5298 13625 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 5212 13625 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 5126 13625 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 5040 13625 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 4954 13625 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 4868 13625 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13585 4782 13625 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 39541 13616 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 39460 13616 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 39379 13616 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 39298 13616 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 39217 13616 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 39136 13616 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 39055 13616 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38974 13616 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38893 13616 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38812 13616 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38731 13616 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38650 13616 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38569 13616 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38488 13616 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38407 13616 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38326 13616 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38245 13616 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38164 13616 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38083 13616 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 38002 13616 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37921 13616 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37840 13616 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37759 13616 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37678 13616 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37597 13616 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37516 13616 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37435 13616 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37354 13616 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37273 13616 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37192 13616 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37111 13616 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 37030 13616 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36949 13616 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36868 13616 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36787 13616 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36706 13616 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36625 13616 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36544 13616 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36463 13616 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36382 13616 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36301 13616 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36220 13616 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36140 13616 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 36060 13616 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35980 13616 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35900 13616 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35820 13616 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35740 13616 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35660 13616 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35580 13616 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35500 13616 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35420 13616 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35340 13616 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35260 13616 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35180 13616 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35100 13616 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 35020 13616 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 34940 13616 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 34860 13616 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13576 34780 13616 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 5642 13544 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 5556 13544 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 5470 13544 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 5384 13544 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 5298 13544 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 5212 13544 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 5126 13544 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 5040 13544 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 4954 13544 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 4868 13544 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13504 4782 13544 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 39541 13534 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 39460 13534 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 39379 13534 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 39298 13534 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 39217 13534 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 39136 13534 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 39055 13534 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38974 13534 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38893 13534 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38812 13534 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38731 13534 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38650 13534 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38569 13534 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38488 13534 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38407 13534 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38326 13534 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38245 13534 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38164 13534 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38083 13534 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 38002 13534 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37921 13534 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37840 13534 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37759 13534 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37678 13534 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37597 13534 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37516 13534 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37435 13534 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37354 13534 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37273 13534 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37192 13534 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37111 13534 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 37030 13534 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36949 13534 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36868 13534 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36787 13534 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36706 13534 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36625 13534 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36544 13534 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36463 13534 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36382 13534 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36301 13534 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36220 13534 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36140 13534 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 36060 13534 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35980 13534 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35900 13534 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35820 13534 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35740 13534 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35660 13534 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35580 13534 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35500 13534 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35420 13534 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35340 13534 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35260 13534 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35180 13534 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35100 13534 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 35020 13534 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 34940 13534 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 34860 13534 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13494 34780 13534 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 5642 13463 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 5556 13463 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 5470 13463 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 5384 13463 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 5298 13463 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 5212 13463 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 5126 13463 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 5040 13463 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 4954 13463 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 4868 13463 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13423 4782 13463 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 39541 13452 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 39460 13452 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 39379 13452 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 39298 13452 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 39217 13452 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 39136 13452 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 39055 13452 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38974 13452 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38893 13452 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38812 13452 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38731 13452 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38650 13452 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38569 13452 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38488 13452 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38407 13452 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38326 13452 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38245 13452 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38164 13452 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38083 13452 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 38002 13452 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37921 13452 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37840 13452 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37759 13452 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37678 13452 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37597 13452 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37516 13452 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37435 13452 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37354 13452 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37273 13452 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37192 13452 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37111 13452 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 37030 13452 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36949 13452 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36868 13452 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36787 13452 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36706 13452 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36625 13452 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36544 13452 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36463 13452 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36382 13452 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36301 13452 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36220 13452 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36140 13452 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 36060 13452 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35980 13452 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35900 13452 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35820 13452 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35740 13452 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35660 13452 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35580 13452 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35500 13452 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35420 13452 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35340 13452 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35260 13452 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35180 13452 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35100 13452 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 35020 13452 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 34940 13452 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 34860 13452 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13412 34780 13452 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 5642 13382 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 5556 13382 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 5470 13382 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 5384 13382 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 5298 13382 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 5212 13382 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 5126 13382 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 5040 13382 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 4954 13382 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 4868 13382 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13342 4782 13382 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 39541 13370 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 39460 13370 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 39379 13370 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 39298 13370 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 39217 13370 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 39136 13370 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 39055 13370 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38974 13370 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38893 13370 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38812 13370 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38731 13370 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38650 13370 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38569 13370 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38488 13370 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38407 13370 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38326 13370 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38245 13370 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38164 13370 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38083 13370 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 38002 13370 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37921 13370 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37840 13370 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37759 13370 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37678 13370 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37597 13370 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37516 13370 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37435 13370 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37354 13370 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37273 13370 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37192 13370 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37111 13370 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 37030 13370 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36949 13370 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36868 13370 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36787 13370 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36706 13370 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36625 13370 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36544 13370 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36463 13370 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36382 13370 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36301 13370 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36220 13370 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36140 13370 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 36060 13370 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35980 13370 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35900 13370 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35820 13370 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35740 13370 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35660 13370 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35580 13370 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35500 13370 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35420 13370 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35340 13370 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35260 13370 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35180 13370 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35100 13370 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 35020 13370 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 34940 13370 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 34860 13370 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13330 34780 13370 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 5642 13301 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 5556 13301 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 5470 13301 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 5384 13301 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 5298 13301 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 5212 13301 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 5126 13301 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 5040 13301 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 4954 13301 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 4868 13301 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13261 4782 13301 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 39541 13288 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 39460 13288 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 39379 13288 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 39298 13288 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 39217 13288 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 39136 13288 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 39055 13288 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38974 13288 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38893 13288 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38812 13288 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38731 13288 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38650 13288 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38569 13288 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38488 13288 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38407 13288 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38326 13288 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38245 13288 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38164 13288 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38083 13288 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 38002 13288 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37921 13288 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37840 13288 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37759 13288 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37678 13288 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37597 13288 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37516 13288 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37435 13288 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37354 13288 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37273 13288 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37192 13288 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37111 13288 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 37030 13288 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36949 13288 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36868 13288 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36787 13288 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36706 13288 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36625 13288 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36544 13288 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36463 13288 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36382 13288 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36301 13288 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36220 13288 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36140 13288 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 36060 13288 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35980 13288 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35900 13288 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35820 13288 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35740 13288 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35660 13288 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35580 13288 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35500 13288 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35420 13288 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35340 13288 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35260 13288 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35180 13288 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35100 13288 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 35020 13288 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 34940 13288 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 34860 13288 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13248 34780 13288 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 5642 13220 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 5556 13220 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 5470 13220 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 5384 13220 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 5298 13220 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 5212 13220 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 5126 13220 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 5040 13220 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 4954 13220 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 4868 13220 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13180 4782 13220 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 39541 13206 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 39460 13206 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 39379 13206 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 39298 13206 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 39217 13206 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 39136 13206 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 39055 13206 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38974 13206 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38893 13206 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38812 13206 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38731 13206 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38650 13206 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38569 13206 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38488 13206 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38407 13206 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38326 13206 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38245 13206 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38164 13206 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38083 13206 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 38002 13206 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37921 13206 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37840 13206 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37759 13206 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37678 13206 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37597 13206 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37516 13206 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37435 13206 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37354 13206 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37273 13206 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37192 13206 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37111 13206 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 37030 13206 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36949 13206 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36868 13206 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36787 13206 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36706 13206 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36625 13206 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36544 13206 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36463 13206 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36382 13206 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36301 13206 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36220 13206 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36140 13206 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 36060 13206 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35980 13206 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35900 13206 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35820 13206 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35740 13206 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35660 13206 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35580 13206 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35500 13206 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35420 13206 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35340 13206 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35260 13206 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35180 13206 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35100 13206 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 35020 13206 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 34940 13206 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 34860 13206 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13166 34780 13206 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 5642 13139 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 5556 13139 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 5470 13139 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 5384 13139 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 5298 13139 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 5212 13139 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 5126 13139 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 5040 13139 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 4954 13139 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 4868 13139 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13099 4782 13139 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 39541 13124 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 39460 13124 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 39379 13124 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 39298 13124 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 39217 13124 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 39136 13124 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 39055 13124 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38974 13124 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38893 13124 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38812 13124 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38731 13124 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38650 13124 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38569 13124 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38488 13124 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38407 13124 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38326 13124 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38245 13124 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38164 13124 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38083 13124 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 38002 13124 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37921 13124 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37840 13124 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37759 13124 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37678 13124 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37597 13124 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37516 13124 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37435 13124 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37354 13124 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37273 13124 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37192 13124 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37111 13124 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 37030 13124 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36949 13124 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36868 13124 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36787 13124 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36706 13124 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36625 13124 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36544 13124 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36463 13124 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36382 13124 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36301 13124 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36220 13124 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36140 13124 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 36060 13124 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35980 13124 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35900 13124 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35820 13124 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35740 13124 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35660 13124 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35580 13124 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35500 13124 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35420 13124 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35340 13124 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35260 13124 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35180 13124 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35100 13124 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 35020 13124 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 34940 13124 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 34860 13124 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13084 34780 13124 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 5642 13058 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 5556 13058 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 5470 13058 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 5384 13058 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 5298 13058 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 5212 13058 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 5126 13058 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 5040 13058 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 4954 13058 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 4868 13058 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13018 4782 13058 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 39541 13042 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 39460 13042 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 39379 13042 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 39298 13042 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 39217 13042 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 39136 13042 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 39055 13042 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38974 13042 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38893 13042 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38812 13042 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38731 13042 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38650 13042 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38569 13042 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38488 13042 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38407 13042 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38326 13042 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38245 13042 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38164 13042 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38083 13042 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 38002 13042 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37921 13042 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37840 13042 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37759 13042 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37678 13042 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37597 13042 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37516 13042 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37435 13042 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37354 13042 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37273 13042 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37192 13042 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37111 13042 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 37030 13042 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36949 13042 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36868 13042 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36787 13042 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36706 13042 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36625 13042 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36544 13042 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36463 13042 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36382 13042 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36301 13042 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36220 13042 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36140 13042 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 36060 13042 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35980 13042 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35900 13042 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35820 13042 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35740 13042 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35660 13042 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35580 13042 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35500 13042 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35420 13042 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35340 13042 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35260 13042 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35180 13042 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35100 13042 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 35020 13042 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 34940 13042 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 34860 13042 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 13002 34780 13042 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 5642 12977 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 5556 12977 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 5470 12977 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 5384 12977 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 5298 12977 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 5212 12977 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 5126 12977 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 5040 12977 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 4954 12977 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 4868 12977 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12937 4782 12977 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 39541 12960 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 39460 12960 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 39379 12960 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 39298 12960 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 39217 12960 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 39136 12960 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 39055 12960 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38974 12960 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38893 12960 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38812 12960 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38731 12960 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38650 12960 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38569 12960 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38488 12960 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38407 12960 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38326 12960 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38245 12960 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38164 12960 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38083 12960 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 38002 12960 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37921 12960 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37840 12960 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37759 12960 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37678 12960 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37597 12960 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37516 12960 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37435 12960 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37354 12960 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37273 12960 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37192 12960 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37111 12960 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 37030 12960 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36949 12960 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36868 12960 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36787 12960 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36706 12960 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36625 12960 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36544 12960 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36463 12960 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36382 12960 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36301 12960 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36220 12960 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36140 12960 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 36060 12960 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35980 12960 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35900 12960 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35820 12960 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35740 12960 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35660 12960 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35580 12960 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35500 12960 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35420 12960 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35340 12960 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35260 12960 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35180 12960 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35100 12960 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 35020 12960 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 34940 12960 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 34860 12960 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12920 34780 12960 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 5642 12896 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 5556 12896 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 5470 12896 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 5384 12896 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 5298 12896 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 5212 12896 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 5126 12896 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 5040 12896 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 4954 12896 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 4868 12896 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12856 4782 12896 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 39541 12878 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 39460 12878 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 39379 12878 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 39298 12878 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 39217 12878 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 39136 12878 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 39055 12878 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38974 12878 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38893 12878 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38812 12878 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38731 12878 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38650 12878 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38569 12878 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38488 12878 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38407 12878 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38326 12878 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38245 12878 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38164 12878 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38083 12878 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 38002 12878 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37921 12878 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37840 12878 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37759 12878 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37678 12878 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37597 12878 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37516 12878 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37435 12878 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37354 12878 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37273 12878 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37192 12878 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37111 12878 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 37030 12878 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36949 12878 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36868 12878 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36787 12878 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36706 12878 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36625 12878 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36544 12878 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36463 12878 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36382 12878 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36301 12878 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36220 12878 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36140 12878 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 36060 12878 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35980 12878 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35900 12878 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35820 12878 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35740 12878 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35660 12878 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35580 12878 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35500 12878 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35420 12878 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35340 12878 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35260 12878 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35180 12878 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35100 12878 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 35020 12878 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 34940 12878 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 34860 12878 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12838 34780 12878 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 5642 12815 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 5556 12815 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 5470 12815 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 5384 12815 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 5298 12815 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 5212 12815 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 5126 12815 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 5040 12815 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 4954 12815 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 4868 12815 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12775 4782 12815 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 39541 12796 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 39460 12796 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 39379 12796 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 39298 12796 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 39217 12796 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 39136 12796 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 39055 12796 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38974 12796 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38893 12796 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38812 12796 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38731 12796 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38650 12796 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38569 12796 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38488 12796 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38407 12796 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38326 12796 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38245 12796 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38164 12796 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38083 12796 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 38002 12796 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37921 12796 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37840 12796 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37759 12796 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37678 12796 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37597 12796 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37516 12796 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37435 12796 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37354 12796 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37273 12796 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37192 12796 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37111 12796 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 37030 12796 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36949 12796 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36868 12796 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36787 12796 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36706 12796 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36625 12796 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36544 12796 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36463 12796 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36382 12796 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36301 12796 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36220 12796 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36140 12796 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 36060 12796 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35980 12796 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35900 12796 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35820 12796 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35740 12796 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35660 12796 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35580 12796 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35500 12796 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35420 12796 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35340 12796 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35260 12796 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35180 12796 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35100 12796 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 35020 12796 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 34940 12796 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 34860 12796 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12756 34780 12796 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 5642 12734 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 5556 12734 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 5470 12734 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 5384 12734 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 5298 12734 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 5212 12734 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 5126 12734 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 5040 12734 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 4954 12734 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 4868 12734 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12694 4782 12734 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 39541 12714 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 39460 12714 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 39379 12714 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 39298 12714 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 39217 12714 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 39136 12714 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 39055 12714 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38974 12714 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38893 12714 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38812 12714 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38731 12714 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38650 12714 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38569 12714 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38488 12714 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38407 12714 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38326 12714 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38245 12714 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38164 12714 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38083 12714 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 38002 12714 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37921 12714 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37840 12714 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37759 12714 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37678 12714 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37597 12714 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37516 12714 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37435 12714 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37354 12714 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37273 12714 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37192 12714 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37111 12714 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 37030 12714 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36949 12714 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36868 12714 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36787 12714 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36706 12714 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36625 12714 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36544 12714 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36463 12714 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36382 12714 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36301 12714 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36220 12714 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36140 12714 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 36060 12714 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35980 12714 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35900 12714 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35820 12714 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35740 12714 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35660 12714 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35580 12714 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35500 12714 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35420 12714 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35340 12714 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35260 12714 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35180 12714 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35100 12714 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 35020 12714 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 34940 12714 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 34860 12714 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12674 34780 12714 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 5642 12653 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 5556 12653 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 5470 12653 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 5384 12653 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 5298 12653 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 5212 12653 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 5126 12653 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 5040 12653 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 4954 12653 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 4868 12653 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12613 4782 12653 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 39541 12632 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 39460 12632 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 39379 12632 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 39298 12632 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 39217 12632 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 39136 12632 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 39055 12632 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38974 12632 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38893 12632 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38812 12632 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38731 12632 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38650 12632 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38569 12632 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38488 12632 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38407 12632 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38326 12632 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38245 12632 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38164 12632 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38083 12632 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 38002 12632 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37921 12632 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37840 12632 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37759 12632 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37678 12632 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37597 12632 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37516 12632 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37435 12632 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37354 12632 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37273 12632 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37192 12632 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37111 12632 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 37030 12632 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36949 12632 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36868 12632 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36787 12632 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36706 12632 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36625 12632 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36544 12632 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36463 12632 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36382 12632 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36301 12632 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36220 12632 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36140 12632 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 36060 12632 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35980 12632 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35900 12632 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35820 12632 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35740 12632 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35660 12632 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35580 12632 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35500 12632 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35420 12632 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35340 12632 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35260 12632 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35180 12632 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35100 12632 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 35020 12632 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 34940 12632 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 34860 12632 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12592 34780 12632 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 5642 12572 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 5556 12572 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 5470 12572 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 5384 12572 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 5298 12572 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 5212 12572 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 5126 12572 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 5040 12572 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 4954 12572 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 4868 12572 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12532 4782 12572 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 39541 12550 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 39460 12550 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 39379 12550 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 39298 12550 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 39217 12550 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 39136 12550 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 39055 12550 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38974 12550 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38893 12550 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38812 12550 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38731 12550 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38650 12550 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38569 12550 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38488 12550 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38407 12550 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38326 12550 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38245 12550 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38164 12550 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38083 12550 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 38002 12550 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37921 12550 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37840 12550 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37759 12550 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37678 12550 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37597 12550 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37516 12550 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37435 12550 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37354 12550 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37273 12550 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37192 12550 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37111 12550 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 37030 12550 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36949 12550 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36868 12550 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36787 12550 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36706 12550 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36625 12550 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36544 12550 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36463 12550 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36382 12550 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36301 12550 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36220 12550 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36140 12550 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 36060 12550 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35980 12550 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35900 12550 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35820 12550 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35740 12550 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35660 12550 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35580 12550 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35500 12550 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35420 12550 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35340 12550 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35260 12550 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35180 12550 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35100 12550 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 35020 12550 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 34940 12550 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 34860 12550 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12510 34780 12550 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 5642 12491 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 5556 12491 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 5470 12491 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 5384 12491 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 5298 12491 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 5212 12491 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 5126 12491 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 5040 12491 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 4954 12491 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 4868 12491 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12451 4782 12491 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 39541 12468 39581 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 39460 12468 39500 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 39379 12468 39419 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 39298 12468 39338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 39217 12468 39257 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 39136 12468 39176 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 39055 12468 39095 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38974 12468 39014 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38893 12468 38933 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38812 12468 38852 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38731 12468 38771 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38650 12468 38690 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38569 12468 38609 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38488 12468 38528 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38407 12468 38447 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38326 12468 38366 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38245 12468 38285 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38164 12468 38204 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38083 12468 38123 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 38002 12468 38042 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37921 12468 37961 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37840 12468 37880 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37759 12468 37799 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37678 12468 37718 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37597 12468 37637 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37516 12468 37556 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37435 12468 37475 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37354 12468 37394 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37273 12468 37313 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37192 12468 37232 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37111 12468 37151 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 37030 12468 37070 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36949 12468 36989 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36868 12468 36908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36787 12468 36827 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36706 12468 36746 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36625 12468 36665 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36544 12468 36584 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36463 12468 36503 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36382 12468 36422 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36301 12468 36341 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36220 12468 36260 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36140 12468 36180 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 36060 12468 36100 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35980 12468 36020 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35900 12468 35940 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35820 12468 35860 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35740 12468 35780 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35660 12468 35700 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35580 12468 35620 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35500 12468 35540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35420 12468 35460 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35340 12468 35380 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35260 12468 35300 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35180 12468 35220 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35100 12468 35140 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 35020 12468 35060 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 34940 12468 34980 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 34860 12468 34900 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12428 34780 12468 34820 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 5642 12410 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 5556 12410 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 5470 12410 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 5384 12410 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 5298 12410 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 5212 12410 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 5126 12410 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 5040 12410 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 4954 12410 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 4868 12410 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12370 4782 12410 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 5642 12329 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 5556 12329 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 5470 12329 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 5384 12329 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 5298 12329 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 5212 12329 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 5126 12329 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 5040 12329 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 4954 12329 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 4868 12329 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12289 4782 12329 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 5642 12248 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 5556 12248 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 5470 12248 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 5384 12248 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 5298 12248 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 5212 12248 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 5126 12248 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 5040 12248 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 4954 12248 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 4868 12248 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12208 4782 12248 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 5642 12167 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 5556 12167 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 5470 12167 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 5384 12167 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 5298 12167 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 5212 12167 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 5126 12167 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 5040 12167 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 4954 12167 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 4868 12167 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12127 4782 12167 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 5642 12086 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 5556 12086 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 5470 12086 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 5384 12086 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 5298 12086 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 5212 12086 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 5126 12086 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 5040 12086 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 4954 12086 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 4868 12086 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 12046 4782 12086 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 5642 12005 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 5556 12005 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 5470 12005 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 5384 12005 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 5298 12005 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 5212 12005 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 5126 12005 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 5040 12005 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 4954 12005 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 4868 12005 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11965 4782 12005 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 5642 11924 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 5556 11924 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 5470 11924 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 5384 11924 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 5298 11924 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 5212 11924 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 5126 11924 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 5040 11924 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 4954 11924 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 4868 11924 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11884 4782 11924 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 5642 11843 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 5556 11843 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 5470 11843 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 5384 11843 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 5298 11843 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 5212 11843 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 5126 11843 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 5040 11843 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 4954 11843 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 4868 11843 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11803 4782 11843 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 5642 11762 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 5556 11762 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 5470 11762 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 5384 11762 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 5298 11762 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 5212 11762 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 5126 11762 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 5040 11762 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 4954 11762 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 4868 11762 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11722 4782 11762 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 5642 11681 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 5556 11681 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 5470 11681 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 5384 11681 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 5298 11681 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 5212 11681 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 5126 11681 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 5040 11681 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 4954 11681 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 4868 11681 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11641 4782 11681 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 5642 11600 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 5556 11600 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 5470 11600 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 5384 11600 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 5298 11600 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 5212 11600 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 5126 11600 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 5040 11600 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 4954 11600 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 4868 11600 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11560 4782 11600 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 5642 11519 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 5556 11519 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 5470 11519 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 5384 11519 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 5298 11519 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 5212 11519 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 5126 11519 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 5040 11519 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 4954 11519 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 4868 11519 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11479 4782 11519 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 5642 11438 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 5556 11438 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 5470 11438 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 5384 11438 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 5298 11438 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 5212 11438 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 5126 11438 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 5040 11438 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 4954 11438 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 4868 11438 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11398 4782 11438 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 5642 11357 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 5556 11357 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 5470 11357 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 5384 11357 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 5298 11357 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 5212 11357 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 5126 11357 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 5040 11357 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 4954 11357 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 4868 11357 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11317 4782 11357 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 5642 11275 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 5556 11275 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 5470 11275 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 5384 11275 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 5298 11275 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 5212 11275 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 5126 11275 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 5040 11275 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 4954 11275 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 4868 11275 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11235 4782 11275 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 5642 11193 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 5556 11193 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 5470 11193 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 5384 11193 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 5298 11193 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 5212 11193 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 5126 11193 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 5040 11193 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 4954 11193 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 4868 11193 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11153 4782 11193 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 5642 11111 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 5556 11111 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 5470 11111 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 5384 11111 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 5298 11111 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 5212 11111 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 5126 11111 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 5040 11111 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 4954 11111 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 4868 11111 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 11071 4782 11111 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 5642 11029 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 5556 11029 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 5470 11029 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 5384 11029 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 5298 11029 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 5212 11029 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 5126 11029 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 5040 11029 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 4954 11029 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 4868 11029 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10989 4782 11029 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 5642 10947 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 5556 10947 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 5470 10947 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 5384 10947 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 5298 10947 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 5212 10947 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 5126 10947 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 5040 10947 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 4954 10947 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 4868 10947 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10907 4782 10947 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 5642 10865 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 5556 10865 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 5470 10865 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 5384 10865 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 5298 10865 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 5212 10865 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 5126 10865 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 5040 10865 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 4954 10865 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 4868 10865 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10825 4782 10865 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 5642 10783 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 5556 10783 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 5470 10783 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 5384 10783 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 5298 10783 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 5212 10783 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 5126 10783 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 5040 10783 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 4954 10783 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 4868 10783 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10743 4782 10783 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 5642 10701 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 5556 10701 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 5470 10701 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 5384 10701 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 5298 10701 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 5212 10701 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 5126 10701 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 5040 10701 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 4954 10701 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 4868 10701 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10661 4782 10701 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 5642 10619 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 5556 10619 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 5470 10619 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 5384 10619 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 5298 10619 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 5212 10619 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 5126 10619 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 5040 10619 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 4954 10619 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 4868 10619 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10579 4782 10619 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 5642 10537 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 5556 10537 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 5470 10537 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 5384 10537 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 5298 10537 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 5212 10537 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 5126 10537 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 5040 10537 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 4954 10537 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 4868 10537 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10497 4782 10537 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 5642 10455 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 5556 10455 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 5470 10455 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 5384 10455 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 5298 10455 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 5212 10455 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 5126 10455 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 5040 10455 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 4954 10455 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 4868 10455 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10415 4782 10455 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 5642 10373 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 5556 10373 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 5470 10373 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 5384 10373 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 5298 10373 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 5212 10373 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 5126 10373 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 5040 10373 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 4954 10373 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 4868 10373 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10333 4782 10373 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 5642 10291 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 5556 10291 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 5470 10291 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 5384 10291 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 5298 10291 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 5212 10291 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 5126 10291 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 5040 10291 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 4954 10291 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 4868 10291 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10251 4782 10291 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 5642 10209 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 5556 10209 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 5470 10209 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 5384 10209 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 5298 10209 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 5212 10209 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 5126 10209 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 5040 10209 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 4954 10209 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 4868 10209 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 10169 4782 10209 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 5642 4862 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 5556 4862 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 5470 4862 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 5384 4862 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 5298 4862 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 5212 4862 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 5126 4862 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 5040 4862 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 4954 4862 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 4868 4862 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4822 4782 4862 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 5642 4781 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 5556 4781 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 5470 4781 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 5384 4781 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 5298 4781 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 5212 4781 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 5126 4781 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 5040 4781 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 4954 4781 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 4868 4781 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4741 4782 4781 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 5642 4700 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 5556 4700 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 5470 4700 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 5384 4700 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 5298 4700 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 5212 4700 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 5126 4700 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 5040 4700 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 4954 4700 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 4868 4700 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4660 4782 4700 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 5642 4619 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 5556 4619 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 5470 4619 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 5384 4619 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 5298 4619 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 5212 4619 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 5126 4619 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 5040 4619 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 4954 4619 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 4868 4619 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4579 4782 4619 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 5642 4538 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 5556 4538 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 5470 4538 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 5384 4538 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 5298 4538 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 5212 4538 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 5126 4538 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 5040 4538 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 4954 4538 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 4868 4538 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4498 4782 4538 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 5642 4457 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 5556 4457 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 5470 4457 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 5384 4457 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 5298 4457 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 5212 4457 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 5126 4457 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 5040 4457 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 4954 4457 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 4868 4457 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4417 4782 4457 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 5642 4376 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 5556 4376 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 5470 4376 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 5384 4376 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 5298 4376 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 5212 4376 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 5126 4376 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 5040 4376 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 4954 4376 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 4868 4376 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4336 4782 4376 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 5642 4295 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 5556 4295 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 5470 4295 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 5384 4295 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 5298 4295 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 5212 4295 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 5126 4295 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 5040 4295 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 4954 4295 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 4868 4295 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4255 4782 4295 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 5642 4214 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 5556 4214 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 5470 4214 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 5384 4214 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 5298 4214 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 5212 4214 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 5126 4214 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 5040 4214 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 4954 4214 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 4868 4214 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4174 4782 4214 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 5642 4133 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 5556 4133 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 5470 4133 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 5384 4133 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 5298 4133 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 5212 4133 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 5126 4133 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 5040 4133 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 4954 4133 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 4868 4133 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4093 4782 4133 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 5642 4052 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 5556 4052 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 5470 4052 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 5384 4052 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 5298 4052 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 5212 4052 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 5126 4052 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 5040 4052 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 4954 4052 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 4868 4052 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 4012 4782 4052 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 5642 3971 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 5556 3971 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 5470 3971 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 5384 3971 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 5298 3971 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 5212 3971 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 5126 3971 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 5040 3971 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 4954 3971 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 4868 3971 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3931 4782 3971 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 5642 3890 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 5556 3890 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 5470 3890 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 5384 3890 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 5298 3890 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 5212 3890 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 5126 3890 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 5040 3890 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 4954 3890 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 4868 3890 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3850 4782 3890 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 5642 3809 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 5556 3809 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 5470 3809 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 5384 3809 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 5298 3809 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 5212 3809 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 5126 3809 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 5040 3809 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 4954 3809 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 4868 3809 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3769 4782 3809 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 5642 3728 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 5556 3728 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 5470 3728 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 5384 3728 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 5298 3728 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 5212 3728 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 5126 3728 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 5040 3728 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 4954 3728 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 4868 3728 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3688 4782 3728 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 5642 3647 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 5556 3647 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 5470 3647 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 5384 3647 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 5298 3647 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 5212 3647 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 5126 3647 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 5040 3647 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 4954 3647 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 4868 3647 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3607 4782 3647 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 5642 3566 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 5556 3566 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 5470 3566 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 5384 3566 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 5298 3566 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 5212 3566 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 5126 3566 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 5040 3566 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 4954 3566 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 4868 3566 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3526 4782 3566 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 5642 3485 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 5556 3485 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 5470 3485 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 5384 3485 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 5298 3485 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 5212 3485 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 5126 3485 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 5040 3485 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 4954 3485 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 4868 3485 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3445 4782 3485 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 5642 3404 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 5556 3404 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 5470 3404 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 5384 3404 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 5298 3404 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 5212 3404 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 5126 3404 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 5040 3404 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 4954 3404 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 4868 3404 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3364 4782 3404 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 5642 3323 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 5556 3323 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 5470 3323 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 5384 3323 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 5298 3323 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 5212 3323 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 5126 3323 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 5040 3323 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 4954 3323 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 4868 3323 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3283 4782 3323 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 5642 3242 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 5556 3242 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 5470 3242 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 5384 3242 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 5298 3242 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 5212 3242 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 5126 3242 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 5040 3242 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 4954 3242 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 4868 3242 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3202 4782 3242 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 5642 3161 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 5556 3161 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 5470 3161 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 5384 3161 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 5298 3161 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 5212 3161 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 5126 3161 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 5040 3161 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 4954 3161 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 4868 3161 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3121 4782 3161 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 5642 3080 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 5556 3080 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 5470 3080 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 5384 3080 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 5298 3080 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 5212 3080 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 5126 3080 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 5040 3080 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 4954 3080 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 4868 3080 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 3040 4782 3080 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 5642 2999 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 5556 2999 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 5470 2999 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 5384 2999 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 5298 2999 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 5212 2999 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 5126 2999 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 5040 2999 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 4954 2999 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 4868 2999 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2959 4782 2999 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 5642 2918 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 5556 2918 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 5470 2918 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 5384 2918 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 5298 2918 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 5212 2918 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 5126 2918 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 5040 2918 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 4954 2918 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 4868 2918 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2878 4782 2918 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 5642 2837 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 5556 2837 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 5470 2837 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 5384 2837 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 5298 2837 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 5212 2837 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 5126 2837 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 5040 2837 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 4954 2837 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 4868 2837 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2797 4782 2837 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 5642 2756 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 5556 2756 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 5470 2756 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 5384 2756 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 5298 2756 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 5212 2756 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 5126 2756 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 5040 2756 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 4954 2756 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 4868 2756 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2716 4782 2756 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 5642 2675 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 5556 2675 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 5470 2675 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 5384 2675 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 5298 2675 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 5212 2675 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 5126 2675 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 5040 2675 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 4954 2675 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 4868 2675 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2635 4782 2675 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 5642 2594 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 5556 2594 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 5470 2594 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 5384 2594 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 5298 2594 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 5212 2594 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 5126 2594 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 5040 2594 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 4954 2594 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 4868 2594 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2554 4782 2594 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 39529 2575 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 39448 2575 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 39367 2575 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 39286 2575 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 39205 2575 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 39124 2575 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 39043 2575 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38962 2575 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38881 2575 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38800 2575 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38719 2575 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38638 2575 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38557 2575 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38476 2575 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38395 2575 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38314 2575 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38233 2575 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38152 2575 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 38071 2575 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37990 2575 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37909 2575 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37828 2575 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37747 2575 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37666 2575 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37585 2575 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37504 2575 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37423 2575 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37342 2575 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37261 2575 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37180 2575 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37099 2575 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 37018 2575 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36937 2575 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36856 2575 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36775 2575 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36694 2575 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36613 2575 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36532 2575 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36451 2575 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36370 2575 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2511 36289 2575 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 34768 2575 36272 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 5642 2513 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 5556 2513 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 5470 2513 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 5384 2513 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 5298 2513 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 5212 2513 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 5126 2513 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 5040 2513 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 4954 2513 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 4868 2513 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2473 4782 2513 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 39529 2495 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 39448 2495 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 39367 2495 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 39286 2495 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 39205 2495 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 39124 2495 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 39043 2495 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38962 2495 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38881 2495 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38800 2495 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38719 2495 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38638 2495 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38557 2495 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38476 2495 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38395 2495 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38314 2495 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38233 2495 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38152 2495 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 38071 2495 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37990 2495 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37909 2495 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37828 2495 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37747 2495 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37666 2495 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37585 2495 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37504 2495 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37423 2495 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37342 2495 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37261 2495 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37180 2495 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37099 2495 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 37018 2495 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36937 2495 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36856 2495 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36775 2495 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36694 2495 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36613 2495 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36532 2495 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36451 2495 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36370 2495 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2431 36289 2495 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 5642 2432 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 5556 2432 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 5470 2432 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 5384 2432 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 5298 2432 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 5212 2432 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 5126 2432 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 5040 2432 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 4954 2432 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 4868 2432 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2392 4782 2432 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 39529 2415 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 39448 2415 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 39367 2415 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 39286 2415 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 39205 2415 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 39124 2415 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 39043 2415 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38962 2415 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38881 2415 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38800 2415 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38719 2415 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38638 2415 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38557 2415 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38476 2415 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38395 2415 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38314 2415 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38233 2415 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38152 2415 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 38071 2415 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37990 2415 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37909 2415 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37828 2415 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37747 2415 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37666 2415 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37585 2415 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37504 2415 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37423 2415 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37342 2415 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37261 2415 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37180 2415 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37099 2415 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 37018 2415 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36937 2415 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36856 2415 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36775 2415 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36694 2415 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36613 2415 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36532 2415 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36451 2415 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36370 2415 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2351 36289 2415 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 5642 2351 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 5556 2351 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 5470 2351 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 5384 2351 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 5298 2351 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 5212 2351 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 5126 2351 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 5040 2351 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 4954 2351 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 4868 2351 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2311 4782 2351 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 39529 2335 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 39448 2335 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 39367 2335 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 39286 2335 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 39205 2335 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 39124 2335 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 39043 2335 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38962 2335 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38881 2335 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38800 2335 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38719 2335 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38638 2335 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38557 2335 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38476 2335 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38395 2335 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38314 2335 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38233 2335 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38152 2335 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 38071 2335 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37990 2335 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37909 2335 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37828 2335 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37747 2335 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37666 2335 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37585 2335 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37504 2335 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37423 2335 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37342 2335 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37261 2335 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37180 2335 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37099 2335 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 37018 2335 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36937 2335 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36856 2335 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36775 2335 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36694 2335 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36613 2335 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36532 2335 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36451 2335 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36370 2335 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2271 36289 2335 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 5642 2270 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 5556 2270 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 5470 2270 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 5384 2270 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 5298 2270 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 5212 2270 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 5126 2270 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 5040 2270 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 4954 2270 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 4868 2270 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2230 4782 2270 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 39529 2255 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 39448 2255 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 39367 2255 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 39286 2255 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 39205 2255 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 39124 2255 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 39043 2255 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38962 2255 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38881 2255 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38800 2255 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38719 2255 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38638 2255 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38557 2255 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38476 2255 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38395 2255 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38314 2255 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38233 2255 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38152 2255 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 38071 2255 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37990 2255 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37909 2255 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37828 2255 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37747 2255 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37666 2255 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37585 2255 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37504 2255 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37423 2255 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37342 2255 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37261 2255 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37180 2255 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37099 2255 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 37018 2255 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36937 2255 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36856 2255 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36775 2255 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36694 2255 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36613 2255 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36532 2255 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36451 2255 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36370 2255 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2191 36289 2255 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 5642 2189 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 5556 2189 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 5470 2189 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 5384 2189 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 5298 2189 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 5212 2189 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 5126 2189 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 5040 2189 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 4954 2189 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 4868 2189 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2149 4782 2189 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 39529 2175 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 39448 2175 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 39367 2175 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 39286 2175 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 39205 2175 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 39124 2175 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 39043 2175 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38962 2175 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38881 2175 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38800 2175 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38719 2175 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38638 2175 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38557 2175 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38476 2175 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38395 2175 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38314 2175 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38233 2175 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38152 2175 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 38071 2175 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37990 2175 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37909 2175 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37828 2175 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37747 2175 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37666 2175 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37585 2175 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37504 2175 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37423 2175 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37342 2175 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37261 2175 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37180 2175 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37099 2175 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 37018 2175 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36937 2175 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36856 2175 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36775 2175 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36694 2175 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36613 2175 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36532 2175 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36451 2175 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36370 2175 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2111 36289 2175 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 5642 2108 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 5556 2108 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 5470 2108 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 5384 2108 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 5298 2108 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 5212 2108 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 5126 2108 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 5040 2108 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 4954 2108 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 4868 2108 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2068 4782 2108 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 39529 2095 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 39448 2095 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 39367 2095 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 39286 2095 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 39205 2095 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 39124 2095 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 39043 2095 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38962 2095 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38881 2095 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38800 2095 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38719 2095 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38638 2095 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38557 2095 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38476 2095 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38395 2095 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38314 2095 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38233 2095 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38152 2095 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 38071 2095 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37990 2095 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37909 2095 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37828 2095 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37747 2095 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37666 2095 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37585 2095 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37504 2095 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37423 2095 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37342 2095 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37261 2095 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37180 2095 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37099 2095 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 37018 2095 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36937 2095 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36856 2095 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36775 2095 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36694 2095 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36613 2095 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36532 2095 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36451 2095 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36370 2095 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 2031 36289 2095 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 5642 2027 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 5556 2027 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 5470 2027 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 5384 2027 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 5298 2027 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 5212 2027 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 5126 2027 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 5040 2027 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 4954 2027 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 4868 2027 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1987 4782 2027 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 39529 2015 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 39448 2015 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 39367 2015 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 39286 2015 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 39205 2015 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 39124 2015 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 39043 2015 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38962 2015 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38881 2015 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38800 2015 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38719 2015 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38638 2015 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38557 2015 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38476 2015 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38395 2015 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38314 2015 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38233 2015 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38152 2015 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 38071 2015 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37990 2015 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37909 2015 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37828 2015 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37747 2015 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37666 2015 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37585 2015 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37504 2015 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37423 2015 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37342 2015 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37261 2015 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37180 2015 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37099 2015 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 37018 2015 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36937 2015 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36856 2015 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36775 2015 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36694 2015 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36613 2015 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36532 2015 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36451 2015 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36370 2015 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1951 36289 2015 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 5642 1946 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 5556 1946 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 5470 1946 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 5384 1946 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 5298 1946 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 5212 1946 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 5126 1946 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 5040 1946 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 4954 1946 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 4868 1946 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1906 4782 1946 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 39529 1935 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 39448 1935 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 39367 1935 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 39286 1935 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 39205 1935 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 39124 1935 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 39043 1935 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38962 1935 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38881 1935 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38800 1935 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38719 1935 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38638 1935 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38557 1935 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38476 1935 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38395 1935 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38314 1935 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38233 1935 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38152 1935 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 38071 1935 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37990 1935 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37909 1935 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37828 1935 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37747 1935 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37666 1935 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37585 1935 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37504 1935 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37423 1935 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37342 1935 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37261 1935 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37180 1935 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37099 1935 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 37018 1935 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36937 1935 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36856 1935 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36775 1935 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36694 1935 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36613 1935 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36532 1935 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36451 1935 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36370 1935 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1871 36289 1935 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 5642 1865 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 5556 1865 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 5470 1865 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 5384 1865 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 5298 1865 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 5212 1865 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 5126 1865 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 5040 1865 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 4954 1865 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 4868 1865 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1825 4782 1865 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 39529 1855 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 39448 1855 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 39367 1855 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 39286 1855 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 39205 1855 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 39124 1855 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 39043 1855 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38962 1855 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38881 1855 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38800 1855 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38719 1855 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38638 1855 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38557 1855 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38476 1855 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38395 1855 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38314 1855 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38233 1855 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38152 1855 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 38071 1855 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37990 1855 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37909 1855 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37828 1855 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37747 1855 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37666 1855 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37585 1855 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37504 1855 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37423 1855 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37342 1855 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37261 1855 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37180 1855 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37099 1855 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 37018 1855 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36937 1855 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36856 1855 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36775 1855 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36694 1855 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36613 1855 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36532 1855 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36451 1855 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36370 1855 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1791 36289 1855 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 5642 1784 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 5556 1784 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 5470 1784 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 5384 1784 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 5298 1784 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 5212 1784 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 5126 1784 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 5040 1784 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 4954 1784 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 4868 1784 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1744 4782 1784 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 39529 1775 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 39448 1775 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 39367 1775 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 39286 1775 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 39205 1775 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 39124 1775 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 39043 1775 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38962 1775 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38881 1775 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38800 1775 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38719 1775 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38638 1775 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38557 1775 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38476 1775 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38395 1775 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38314 1775 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38233 1775 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38152 1775 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 38071 1775 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37990 1775 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37909 1775 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37828 1775 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37747 1775 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37666 1775 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37585 1775 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37504 1775 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37423 1775 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37342 1775 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37261 1775 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37180 1775 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37099 1775 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 37018 1775 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36937 1775 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36856 1775 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36775 1775 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36694 1775 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36613 1775 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36532 1775 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36451 1775 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36370 1775 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1711 36289 1775 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 5642 1703 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 5556 1703 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 5470 1703 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 5384 1703 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 5298 1703 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 5212 1703 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 5126 1703 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 5040 1703 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 4954 1703 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 4868 1703 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1663 4782 1703 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 39529 1695 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 39448 1695 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 39367 1695 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 39286 1695 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 39205 1695 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 39124 1695 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 39043 1695 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38962 1695 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38881 1695 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38800 1695 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38719 1695 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38638 1695 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38557 1695 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38476 1695 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38395 1695 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38314 1695 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38233 1695 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38152 1695 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 38071 1695 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37990 1695 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37909 1695 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37828 1695 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37747 1695 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37666 1695 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37585 1695 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37504 1695 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37423 1695 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37342 1695 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37261 1695 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37180 1695 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37099 1695 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 37018 1695 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36937 1695 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36856 1695 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36775 1695 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36694 1695 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36613 1695 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36532 1695 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36451 1695 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36370 1695 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1631 36289 1695 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 5642 1622 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 5556 1622 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 5470 1622 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 5384 1622 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 5298 1622 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 5212 1622 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 5126 1622 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 5040 1622 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 4954 1622 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 4868 1622 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1582 4782 1622 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 39529 1615 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 39448 1615 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 39367 1615 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 39286 1615 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 39205 1615 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 39124 1615 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 39043 1615 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38962 1615 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38881 1615 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38800 1615 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38719 1615 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38638 1615 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38557 1615 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38476 1615 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38395 1615 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38314 1615 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38233 1615 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38152 1615 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 38071 1615 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37990 1615 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37909 1615 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37828 1615 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37747 1615 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37666 1615 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37585 1615 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37504 1615 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37423 1615 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37342 1615 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37261 1615 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37180 1615 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37099 1615 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 37018 1615 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36937 1615 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36856 1615 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36775 1615 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36694 1615 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36613 1615 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36532 1615 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36451 1615 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36370 1615 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1551 36289 1615 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 5642 1541 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 5556 1541 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 5470 1541 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 5384 1541 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 5298 1541 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 5212 1541 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 5126 1541 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 5040 1541 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 4954 1541 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 4868 1541 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1501 4782 1541 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 39529 1535 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 39448 1535 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 39367 1535 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 39286 1535 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 39205 1535 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 39124 1535 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 39043 1535 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38962 1535 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38881 1535 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38800 1535 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38719 1535 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38638 1535 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38557 1535 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38476 1535 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38395 1535 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38314 1535 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38233 1535 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38152 1535 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 38071 1535 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37990 1535 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37909 1535 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37828 1535 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37747 1535 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37666 1535 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37585 1535 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37504 1535 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37423 1535 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37342 1535 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37261 1535 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37180 1535 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37099 1535 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 37018 1535 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36937 1535 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36856 1535 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36775 1535 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36694 1535 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36613 1535 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36532 1535 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36451 1535 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36370 1535 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1471 36289 1535 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 5642 1460 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 5556 1460 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 5470 1460 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 5384 1460 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 5298 1460 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 5212 1460 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 5126 1460 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 5040 1460 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 4954 1460 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 4868 1460 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1420 4782 1460 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 39529 1455 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 39448 1455 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 39367 1455 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 39286 1455 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 39205 1455 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 39124 1455 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 39043 1455 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38962 1455 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38881 1455 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38800 1455 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38719 1455 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38638 1455 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38557 1455 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38476 1455 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38395 1455 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38314 1455 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38233 1455 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38152 1455 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 38071 1455 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37990 1455 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37909 1455 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37828 1455 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37747 1455 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37666 1455 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37585 1455 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37504 1455 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37423 1455 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37342 1455 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37261 1455 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37180 1455 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37099 1455 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 37018 1455 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36937 1455 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36856 1455 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36775 1455 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36694 1455 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36613 1455 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36532 1455 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36451 1455 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36370 1455 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1391 36289 1455 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 5642 1379 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 5556 1379 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 5470 1379 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 5384 1379 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 5298 1379 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 5212 1379 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 5126 1379 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 5040 1379 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 4954 1379 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 4868 1379 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1339 4782 1379 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 39529 1375 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 39448 1375 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 39367 1375 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 39286 1375 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 39205 1375 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 39124 1375 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 39043 1375 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38962 1375 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38881 1375 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38800 1375 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38719 1375 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38638 1375 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38557 1375 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38476 1375 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38395 1375 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38314 1375 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38233 1375 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38152 1375 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 38071 1375 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37990 1375 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37909 1375 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37828 1375 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37747 1375 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37666 1375 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37585 1375 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37504 1375 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37423 1375 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37342 1375 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37261 1375 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37180 1375 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37099 1375 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 37018 1375 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36937 1375 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36856 1375 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36775 1375 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36694 1375 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36613 1375 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36532 1375 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36451 1375 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36370 1375 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1311 36289 1375 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 5642 1298 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 5556 1298 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 5470 1298 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 5384 1298 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 5298 1298 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 5212 1298 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 5126 1298 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 5040 1298 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 4954 1298 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 4868 1298 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1258 4782 1298 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 39529 1295 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 39448 1295 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 39367 1295 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 39286 1295 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 39205 1295 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 39124 1295 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 39043 1295 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38962 1295 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38881 1295 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38800 1295 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38719 1295 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38638 1295 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38557 1295 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38476 1295 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38395 1295 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38314 1295 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38233 1295 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38152 1295 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 38071 1295 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37990 1295 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37909 1295 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37828 1295 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37747 1295 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37666 1295 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37585 1295 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37504 1295 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37423 1295 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37342 1295 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37261 1295 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37180 1295 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37099 1295 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 37018 1295 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36937 1295 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36856 1295 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36775 1295 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36694 1295 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36613 1295 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36532 1295 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36451 1295 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36370 1295 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1231 36289 1295 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 5642 1217 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 5556 1217 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 5470 1217 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 5384 1217 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 5298 1217 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 5212 1217 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 5126 1217 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 5040 1217 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 4954 1217 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 4868 1217 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1177 4782 1217 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 39529 1215 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 39448 1215 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 39367 1215 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 39286 1215 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 39205 1215 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 39124 1215 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 39043 1215 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38962 1215 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38881 1215 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38800 1215 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38719 1215 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38638 1215 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38557 1215 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38476 1215 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38395 1215 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38314 1215 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38233 1215 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38152 1215 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 38071 1215 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37990 1215 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37909 1215 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37828 1215 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37747 1215 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37666 1215 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37585 1215 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37504 1215 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37423 1215 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37342 1215 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37261 1215 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37180 1215 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37099 1215 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 37018 1215 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36937 1215 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36856 1215 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36775 1215 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36694 1215 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36613 1215 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36532 1215 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36451 1215 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36370 1215 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1151 36289 1215 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 5642 1136 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 5556 1136 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 5470 1136 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 5384 1136 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 5298 1136 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 5212 1136 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 5126 1136 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 5040 1136 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 4954 1136 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 4868 1136 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1096 4782 1136 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 39529 1135 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 39448 1135 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 39367 1135 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 39286 1135 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 39205 1135 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 39124 1135 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 39043 1135 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38962 1135 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38881 1135 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38800 1135 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38719 1135 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38638 1135 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38557 1135 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38476 1135 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38395 1135 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38314 1135 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38233 1135 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38152 1135 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 38071 1135 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37990 1135 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37909 1135 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37828 1135 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37747 1135 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37666 1135 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37585 1135 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37504 1135 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37423 1135 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37342 1135 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37261 1135 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37180 1135 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37099 1135 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 37018 1135 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36937 1135 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36856 1135 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36775 1135 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36694 1135 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36613 1135 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36532 1135 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36451 1135 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36370 1135 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1071 36289 1135 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 5642 1055 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 5556 1055 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 5470 1055 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 5384 1055 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 5298 1055 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 5212 1055 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 5126 1055 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 5040 1055 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 4954 1055 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 4868 1055 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 1015 4782 1055 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 39529 1055 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 39448 1055 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 39367 1055 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 39286 1055 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 39205 1055 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 39124 1055 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 39043 1055 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38962 1055 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38881 1055 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38800 1055 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38719 1055 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38638 1055 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38557 1055 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38476 1055 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38395 1055 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38314 1055 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38233 1055 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38152 1055 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 38071 1055 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37990 1055 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37909 1055 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37828 1055 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37747 1055 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37666 1055 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37585 1055 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37504 1055 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37423 1055 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37342 1055 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37261 1055 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37180 1055 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37099 1055 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 37018 1055 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36937 1055 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36856 1055 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36775 1055 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36694 1055 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36613 1055 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36532 1055 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36451 1055 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36370 1055 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 991 36289 1055 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 5642 974 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 5556 974 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 5470 974 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 5384 974 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 5298 974 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 5212 974 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 5126 974 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 5040 974 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 4954 974 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 4868 974 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 934 4782 974 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 39529 975 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 39448 975 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 39367 975 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 39286 975 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 39205 975 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 39124 975 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 39043 975 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38962 975 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38881 975 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38800 975 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38719 975 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38638 975 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38557 975 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38476 975 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38395 975 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38314 975 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38233 975 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38152 975 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 38071 975 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37990 975 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37909 975 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37828 975 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37747 975 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37666 975 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37585 975 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37504 975 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37423 975 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37342 975 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37261 975 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37180 975 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37099 975 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 37018 975 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36937 975 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36856 975 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36775 975 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36694 975 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36613 975 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36532 975 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36451 975 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36370 975 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 911 36289 975 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 5642 893 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 5556 893 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 5470 893 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 5384 893 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 5298 893 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 5212 893 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 5126 893 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 5040 893 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 4954 893 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 4868 893 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 853 4782 893 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 39529 895 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 39448 895 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 39367 895 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 39286 895 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 39205 895 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 39124 895 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 39043 895 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38962 895 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38881 895 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38800 895 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38719 895 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38638 895 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38557 895 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38476 895 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38395 895 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38314 895 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38233 895 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38152 895 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 38071 895 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37990 895 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37909 895 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37828 895 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37747 895 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37666 895 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37585 895 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37504 895 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37423 895 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37342 895 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37261 895 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37180 895 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37099 895 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 37018 895 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36937 895 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36856 895 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36775 895 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36694 895 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36613 895 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36532 895 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36451 895 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36370 895 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 831 36289 895 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 5642 812 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 5556 812 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 5470 812 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 5384 812 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 5298 812 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 5212 812 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 5126 812 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 5040 812 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 4954 812 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 4868 812 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 772 4782 812 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 39529 815 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 39448 815 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 39367 815 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 39286 815 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 39205 815 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 39124 815 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 39043 815 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38962 815 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38881 815 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38800 815 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38719 815 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38638 815 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38557 815 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38476 815 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38395 815 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38314 815 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38233 815 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38152 815 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 38071 815 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37990 815 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37909 815 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37828 815 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37747 815 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37666 815 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37585 815 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37504 815 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37423 815 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37342 815 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37261 815 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37180 815 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37099 815 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 37018 815 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36937 815 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36856 815 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36775 815 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36694 815 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36613 815 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36532 815 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36451 815 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36370 815 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 751 36289 815 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 5642 731 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 5556 731 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 5470 731 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 5384 731 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 5298 731 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 5212 731 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 5126 731 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 5040 731 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 4954 731 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 4868 731 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 691 4782 731 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 39529 735 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 39448 735 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 39367 735 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 39286 735 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 39205 735 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 39124 735 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 39043 735 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38962 735 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38881 735 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38800 735 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38719 735 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38638 735 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38557 735 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38476 735 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38395 735 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38314 735 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38233 735 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38152 735 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 38071 735 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37990 735 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37909 735 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37828 735 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37747 735 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37666 735 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37585 735 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37504 735 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37423 735 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37342 735 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37261 735 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37180 735 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37099 735 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 37018 735 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36937 735 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36856 735 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36775 735 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36694 735 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36613 735 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36532 735 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36451 735 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36370 735 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 671 36289 735 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 5642 650 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 5556 650 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 5470 650 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 5384 650 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 5298 650 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 5212 650 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 5126 650 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 5040 650 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 4954 650 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 4868 650 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 610 4782 650 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 39529 655 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 39448 655 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 39367 655 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 39286 655 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 39205 655 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 39124 655 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 39043 655 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38962 655 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38881 655 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38800 655 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38719 655 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38638 655 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38557 655 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38476 655 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38395 655 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38314 655 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38233 655 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38152 655 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 38071 655 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37990 655 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37909 655 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37828 655 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37747 655 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37666 655 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37585 655 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37504 655 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37423 655 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37342 655 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37261 655 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37180 655 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37099 655 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 37018 655 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36937 655 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36856 655 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36775 655 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36694 655 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36613 655 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36532 655 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36451 655 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36370 655 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 591 36289 655 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 5642 568 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 5556 568 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 5470 568 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 5384 568 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 5298 568 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 5212 568 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 5126 568 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 5040 568 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 4954 568 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 4868 568 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 528 4782 568 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 39529 575 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 39448 575 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 39367 575 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 39286 575 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 39205 575 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 39124 575 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 39043 575 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38962 575 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38881 575 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38800 575 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38719 575 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38638 575 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38557 575 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38476 575 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38395 575 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38314 575 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38233 575 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38152 575 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 38071 575 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37990 575 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37909 575 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37828 575 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37747 575 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37666 575 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37585 575 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37504 575 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37423 575 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37342 575 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37261 575 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37180 575 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37099 575 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 37018 575 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36937 575 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36856 575 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36775 575 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36694 575 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36613 575 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36532 575 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36451 575 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36370 575 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 511 36289 575 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 5642 486 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 5556 486 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 5470 486 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 5384 486 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 5298 486 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 5212 486 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 5126 486 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 5040 486 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 4954 486 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 4868 486 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 446 4782 486 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 39529 495 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 39448 495 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 39367 495 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 39286 495 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 39205 495 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 39124 495 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 39043 495 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38962 495 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38881 495 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38800 495 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38719 495 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38638 495 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38557 495 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38476 495 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38395 495 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38314 495 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38233 495 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38152 495 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 38071 495 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37990 495 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37909 495 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37828 495 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37747 495 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37666 495 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37585 495 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37504 495 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37423 495 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37342 495 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37261 495 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37180 495 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37099 495 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 37018 495 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36937 495 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36856 495 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36775 495 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36694 495 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36613 495 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36532 495 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36451 495 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36370 495 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 431 36289 495 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 5642 404 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 5556 404 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 5470 404 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 5384 404 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 5298 404 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 5212 404 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 5126 404 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 5040 404 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 4954 404 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 4868 404 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 364 4782 404 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 39529 415 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 39448 415 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 39367 415 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 39286 415 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 39205 415 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 39124 415 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 39043 415 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38962 415 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38881 415 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38800 415 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38719 415 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38638 415 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38557 415 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38476 415 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38395 415 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38314 415 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38233 415 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38152 415 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 38071 415 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37990 415 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37909 415 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37828 415 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37747 415 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37666 415 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37585 415 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37504 415 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37423 415 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37342 415 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37261 415 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37180 415 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37099 415 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 37018 415 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36937 415 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36856 415 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36775 415 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36694 415 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36613 415 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36532 415 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36451 415 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36370 415 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 351 36289 415 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 39529 335 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 39448 335 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 39367 335 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 39286 335 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 39205 335 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 39124 335 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 39043 335 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38962 335 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38881 335 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38800 335 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38719 335 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38638 335 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38557 335 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38476 335 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38395 335 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38314 335 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38233 335 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38152 335 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 38071 335 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37990 335 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37909 335 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37828 335 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37747 335 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37666 335 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37585 335 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37504 335 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37423 335 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37342 335 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37261 335 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37180 335 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37099 335 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 37018 335 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36937 335 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36856 335 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36775 335 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36694 335 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36613 335 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36532 335 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36451 335 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36370 335 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 271 36289 335 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 5642 322 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 5556 322 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 5470 322 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 5384 322 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 5298 322 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 5212 322 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 5126 322 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 5040 322 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 4954 322 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 4868 322 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 282 4782 322 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 39529 255 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 39448 255 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 39367 255 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 39286 255 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 39205 255 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 39124 255 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 39043 255 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38962 255 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38881 255 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38800 255 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38719 255 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38638 255 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38557 255 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38476 255 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38395 255 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38314 255 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38233 255 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38152 255 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 38071 255 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37990 255 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37909 255 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37828 255 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37747 255 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37666 255 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37585 255 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37504 255 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37423 255 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37342 255 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37261 255 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37180 255 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37099 255 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 37018 255 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36937 255 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36856 255 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36775 255 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36694 255 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36613 255 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36532 255 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36451 255 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36370 255 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 191 36289 255 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 5642 240 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 5556 240 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 5470 240 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 5384 240 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 5298 240 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 5212 240 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 5126 240 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 5040 240 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 4954 240 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 4868 240 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 200 4782 240 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 39529 175 39593 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 39448 175 39512 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 39367 175 39431 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 39286 175 39350 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 39205 175 39269 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 39124 175 39188 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 39043 175 39107 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38962 175 39026 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38881 175 38945 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38800 175 38864 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38719 175 38783 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38638 175 38702 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38557 175 38621 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38476 175 38540 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38395 175 38459 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38314 175 38378 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38233 175 38297 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38152 175 38216 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 38071 175 38135 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37990 175 38054 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37909 175 37973 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37828 175 37892 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37747 175 37811 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37666 175 37730 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37585 175 37649 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37504 175 37568 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37423 175 37487 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37342 175 37406 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37261 175 37325 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37180 175 37244 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37099 175 37163 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 37018 175 37082 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36937 175 37001 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36856 175 36920 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36775 175 36839 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36694 175 36758 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36613 175 36677 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36532 175 36596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36451 175 36515 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36370 175 36434 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 111 36289 175 36353 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 5642 158 5682 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 5556 158 5596 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 5470 158 5510 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 5384 158 5424 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 5298 158 5338 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 5212 158 5252 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 5126 158 5166 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 5040 158 5080 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 4954 158 4994 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 4868 158 4908 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal3 s 118 4782 158 4822 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 53 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 54 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10151 11248 14858 12136 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 10156 11247 15000 12137 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 12082 14840 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 12000 14840 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11918 14840 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11836 14840 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11754 14840 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11672 14840 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11590 14840 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11508 14840 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11426 14840 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11344 14840 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14800 11262 14840 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 12082 14759 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 12000 14759 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11918 14759 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11836 14759 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11754 14759 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11672 14759 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11590 14759 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11508 14759 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11426 14759 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11344 14759 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14719 11262 14759 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 12082 14678 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 12000 14678 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11918 14678 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11836 14678 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11754 14678 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11672 14678 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11590 14678 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11508 14678 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11426 14678 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11344 14678 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14638 11262 14678 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 12082 14597 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 12000 14597 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11918 14597 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11836 14597 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11754 14597 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11672 14597 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11590 14597 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11508 14597 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11426 14597 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11344 14597 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14557 11262 14597 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 12082 14516 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 12000 14516 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11918 14516 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11836 14516 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11754 14516 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11672 14516 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11590 14516 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11508 14516 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11426 14516 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11344 14516 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14476 11262 14516 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 12082 14435 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 12000 14435 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11918 14435 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11836 14435 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11754 14435 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11672 14435 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11590 14435 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11508 14435 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11426 14435 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11344 14435 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14395 11262 14435 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 12082 14354 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 12000 14354 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11918 14354 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11836 14354 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11754 14354 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11672 14354 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11590 14354 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11508 14354 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11426 14354 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11344 14354 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14314 11262 14354 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 12082 14273 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 12000 14273 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11918 14273 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11836 14273 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11754 14273 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11672 14273 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11590 14273 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11508 14273 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11426 14273 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11344 14273 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14233 11262 14273 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 12082 14192 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 12000 14192 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11918 14192 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11836 14192 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11754 14192 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11672 14192 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11590 14192 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11508 14192 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11426 14192 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11344 14192 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14152 11262 14192 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 12082 14111 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 12000 14111 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11918 14111 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11836 14111 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11754 14111 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11672 14111 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11590 14111 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11508 14111 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11426 14111 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11344 14111 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 14071 11262 14111 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 12082 14030 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 12000 14030 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11918 14030 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11836 14030 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11754 14030 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11672 14030 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11590 14030 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11508 14030 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11426 14030 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11344 14030 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13990 11262 14030 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 12082 13949 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 12000 13949 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11918 13949 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11836 13949 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11754 13949 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11672 13949 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11590 13949 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11508 13949 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11426 13949 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11344 13949 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13909 11262 13949 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 12082 13868 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 12000 13868 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11918 13868 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11836 13868 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11754 13868 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11672 13868 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11590 13868 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11508 13868 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11426 13868 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11344 13868 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13828 11262 13868 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 12082 13787 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 12000 13787 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11918 13787 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11836 13787 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11754 13787 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11672 13787 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11590 13787 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11508 13787 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11426 13787 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11344 13787 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13747 11262 13787 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 12082 13706 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 12000 13706 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11918 13706 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11836 13706 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11754 13706 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11672 13706 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11590 13706 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11508 13706 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11426 13706 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11344 13706 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13666 11262 13706 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 12082 13625 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 12000 13625 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11918 13625 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11836 13625 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11754 13625 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11672 13625 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11590 13625 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11508 13625 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11426 13625 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11344 13625 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13585 11262 13625 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 12082 13544 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 12000 13544 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11918 13544 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11836 13544 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11754 13544 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11672 13544 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11590 13544 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11508 13544 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11426 13544 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11344 13544 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13504 11262 13544 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 12082 13463 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 12000 13463 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11918 13463 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11836 13463 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11754 13463 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11672 13463 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11590 13463 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11508 13463 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11426 13463 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11344 13463 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13423 11262 13463 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 12082 13382 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 12000 13382 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11918 13382 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11836 13382 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11754 13382 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11672 13382 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11590 13382 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11508 13382 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11426 13382 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11344 13382 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13342 11262 13382 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 12082 13301 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 12000 13301 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11918 13301 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11836 13301 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11754 13301 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11672 13301 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11590 13301 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11508 13301 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11426 13301 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11344 13301 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13261 11262 13301 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 12082 13220 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 12000 13220 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11918 13220 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11836 13220 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11754 13220 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11672 13220 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11590 13220 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11508 13220 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11426 13220 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11344 13220 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13180 11262 13220 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 12082 13139 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 12000 13139 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11918 13139 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11836 13139 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11754 13139 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11672 13139 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11590 13139 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11508 13139 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11426 13139 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11344 13139 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13099 11262 13139 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 12082 13058 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 12000 13058 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11918 13058 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11836 13058 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11754 13058 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11672 13058 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11590 13058 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11508 13058 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11426 13058 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11344 13058 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 13018 11262 13058 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 12082 12977 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 12000 12977 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11918 12977 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11836 12977 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11754 12977 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11672 12977 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11590 12977 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11508 12977 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11426 12977 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11344 12977 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12937 11262 12977 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 12082 12896 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 12000 12896 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11918 12896 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11836 12896 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11754 12896 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11672 12896 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11590 12896 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11508 12896 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11426 12896 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11344 12896 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12856 11262 12896 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 12082 12815 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 12000 12815 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11918 12815 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11836 12815 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11754 12815 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11672 12815 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11590 12815 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11508 12815 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11426 12815 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11344 12815 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12775 11262 12815 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 12082 12734 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 12000 12734 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11918 12734 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11836 12734 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11754 12734 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11672 12734 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11590 12734 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11508 12734 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11426 12734 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11344 12734 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12694 11262 12734 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 12082 12653 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 12000 12653 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11918 12653 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11836 12653 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11754 12653 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11672 12653 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11590 12653 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11508 12653 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11426 12653 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11344 12653 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12613 11262 12653 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 12082 12572 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 12000 12572 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11918 12572 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11836 12572 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11754 12572 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11672 12572 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11590 12572 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11508 12572 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11426 12572 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11344 12572 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12532 11262 12572 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 12082 12491 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 12000 12491 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11918 12491 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11836 12491 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11754 12491 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11672 12491 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11590 12491 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11508 12491 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11426 12491 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11344 12491 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12451 11262 12491 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 12082 12410 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 12000 12410 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11918 12410 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11836 12410 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11754 12410 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11672 12410 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11590 12410 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11508 12410 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11426 12410 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11344 12410 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12370 11262 12410 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 12082 12329 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 12000 12329 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11918 12329 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11836 12329 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11754 12329 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11672 12329 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11590 12329 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11508 12329 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11426 12329 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11344 12329 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12289 11262 12329 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 12082 12248 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 12000 12248 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11918 12248 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11836 12248 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11754 12248 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11672 12248 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11590 12248 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11508 12248 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11426 12248 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11344 12248 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12208 11262 12248 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 12082 12167 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 12000 12167 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11918 12167 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11836 12167 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11754 12167 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11672 12167 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11590 12167 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11508 12167 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11426 12167 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11344 12167 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12127 11262 12167 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 12082 12086 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 12000 12086 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11918 12086 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11836 12086 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11754 12086 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11672 12086 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11590 12086 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11508 12086 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11426 12086 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11344 12086 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 12046 11262 12086 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 12082 12005 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 12000 12005 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11918 12005 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11836 12005 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11754 12005 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11672 12005 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11590 12005 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11508 12005 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11426 12005 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11344 12005 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11965 11262 12005 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 12082 11924 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 12000 11924 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11918 11924 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11836 11924 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11754 11924 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11672 11924 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11590 11924 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11508 11924 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11426 11924 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11344 11924 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11884 11262 11924 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 12082 11843 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 12000 11843 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11918 11843 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11836 11843 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11754 11843 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11672 11843 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11590 11843 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11508 11843 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11426 11843 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11344 11843 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11803 11262 11843 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 12082 11762 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 12000 11762 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11918 11762 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11836 11762 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11754 11762 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11672 11762 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11590 11762 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11508 11762 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11426 11762 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11344 11762 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11722 11262 11762 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 12082 11681 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 12000 11681 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11918 11681 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11836 11681 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11754 11681 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11672 11681 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11590 11681 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11508 11681 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11426 11681 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11344 11681 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11641 11262 11681 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 12082 11600 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 12000 11600 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11918 11600 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11836 11600 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11754 11600 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11672 11600 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11590 11600 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11508 11600 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11426 11600 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11344 11600 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11560 11262 11600 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 12082 11519 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 12000 11519 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11918 11519 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11836 11519 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11754 11519 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11672 11519 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11590 11519 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11508 11519 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11426 11519 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11344 11519 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11479 11262 11519 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 12082 11438 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 12000 11438 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11918 11438 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11836 11438 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11754 11438 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11672 11438 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11590 11438 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11508 11438 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11426 11438 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11344 11438 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11398 11262 11438 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 12082 11357 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 12000 11357 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11918 11357 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11836 11357 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11754 11357 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11672 11357 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11590 11357 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11508 11357 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11426 11357 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11344 11357 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11317 11262 11357 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 12082 11275 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 12000 11275 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11918 11275 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11836 11275 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11754 11275 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11672 11275 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11590 11275 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11508 11275 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11426 11275 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11344 11275 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11235 11262 11275 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 12082 11193 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 12000 11193 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11918 11193 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11836 11193 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11754 11193 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11672 11193 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11590 11193 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11508 11193 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11426 11193 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11344 11193 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11153 11262 11193 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 12082 11111 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 12000 11111 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11918 11111 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11836 11111 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11754 11111 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11672 11111 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11590 11111 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11508 11111 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11426 11111 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11344 11111 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 11071 11262 11111 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 12082 11029 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 12000 11029 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11918 11029 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11836 11029 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11754 11029 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11672 11029 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11590 11029 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11508 11029 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11426 11029 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11344 11029 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10989 11262 11029 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 12082 10947 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 12000 10947 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11918 10947 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11836 10947 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11754 10947 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11672 10947 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11590 10947 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11508 10947 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11426 10947 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11344 10947 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10907 11262 10947 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 12082 10865 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 12000 10865 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11918 10865 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11836 10865 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11754 10865 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11672 10865 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11590 10865 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11508 10865 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11426 10865 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11344 10865 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10825 11262 10865 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 12082 10783 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 12000 10783 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11918 10783 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11836 10783 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11754 10783 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11672 10783 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11590 10783 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11508 10783 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11426 10783 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11344 10783 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10743 11262 10783 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 12082 10701 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 12000 10701 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11918 10701 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11836 10701 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11754 10701 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11672 10701 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11590 10701 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11508 10701 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11426 10701 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11344 10701 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10661 11262 10701 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 12082 10619 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 12000 10619 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11918 10619 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11836 10619 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11754 10619 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11672 10619 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11590 10619 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11508 10619 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11426 10619 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11344 10619 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10579 11262 10619 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 12082 10537 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 12000 10537 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11918 10537 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11836 10537 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11754 10537 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11672 10537 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11590 10537 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11508 10537 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11426 10537 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11344 10537 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10497 11262 10537 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 12082 10455 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 12000 10455 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11918 10455 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11836 10455 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11754 10455 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11672 10455 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11590 10455 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11508 10455 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11426 10455 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11344 10455 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10415 11262 10455 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 12082 10373 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 12000 10373 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11918 10373 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11836 10373 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11754 10373 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11672 10373 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11590 10373 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11508 10373 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11426 10373 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11344 10373 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10333 11262 10373 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 12082 10291 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 12000 10291 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11918 10291 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11836 10291 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11754 10291 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11672 10291 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11590 10291 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11508 10291 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11426 10291 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11344 10291 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10251 11262 10291 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 12082 10209 12122 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 12000 10209 12040 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11918 10209 11958 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11836 10209 11876 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11754 10209 11794 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11672 10209 11712 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11590 10209 11630 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11508 10209 11548 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11426 10209 11466 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11344 10209 11384 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 10169 11262 10209 11302 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 12070 4874 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 12070 4874 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11988 4874 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11988 4874 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11906 4874 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11906 4874 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11824 4874 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11824 4874 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11742 4874 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11742 4874 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11660 4874 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11660 4874 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11578 4874 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11578 4874 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11496 4874 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11496 4874 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11414 4874 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11414 4874 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11332 4874 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11332 4874 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4810 11250 4874 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4810 11250 4874 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 12070 4793 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 12070 4793 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11988 4793 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11988 4793 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11906 4793 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11906 4793 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11824 4793 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11824 4793 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11742 4793 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11742 4793 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11660 4793 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11660 4793 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11578 4793 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11578 4793 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11496 4793 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11496 4793 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11414 4793 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11414 4793 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11332 4793 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11332 4793 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4729 11250 4793 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4729 11250 4793 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 12070 4712 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 12070 4712 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11988 4712 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11988 4712 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11906 4712 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11906 4712 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11824 4712 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11824 4712 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11742 4712 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11742 4712 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11660 4712 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11660 4712 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11578 4712 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11578 4712 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11496 4712 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11496 4712 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11414 4712 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11414 4712 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11332 4712 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11332 4712 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4648 11250 4712 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4648 11250 4712 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 12070 4631 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 12070 4631 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11988 4631 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11988 4631 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11906 4631 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11906 4631 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11824 4631 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11824 4631 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11742 4631 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11742 4631 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11660 4631 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11660 4631 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11578 4631 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11578 4631 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11496 4631 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11496 4631 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11414 4631 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11414 4631 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11332 4631 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11332 4631 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4567 11250 4631 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4567 11250 4631 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 12070 4550 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 12070 4550 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11988 4550 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11988 4550 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11906 4550 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11906 4550 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11824 4550 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11824 4550 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11742 4550 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11742 4550 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11660 4550 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11660 4550 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11578 4550 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11578 4550 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11496 4550 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11496 4550 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11414 4550 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11414 4550 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11332 4550 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11332 4550 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4486 11250 4550 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4486 11250 4550 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 12070 4469 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 12070 4469 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11988 4469 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11988 4469 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11906 4469 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11906 4469 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11824 4469 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11824 4469 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11742 4469 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11742 4469 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11660 4469 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11660 4469 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11578 4469 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11578 4469 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11496 4469 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11496 4469 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11414 4469 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11414 4469 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11332 4469 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11332 4469 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4405 11250 4469 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4405 11250 4469 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 12070 4388 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 12070 4388 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11988 4388 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11988 4388 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11906 4388 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11906 4388 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11824 4388 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11824 4388 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11742 4388 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11742 4388 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11660 4388 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11660 4388 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11578 4388 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11578 4388 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11496 4388 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11496 4388 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11414 4388 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11414 4388 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11332 4388 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11332 4388 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4324 11250 4388 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4324 11250 4388 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 12070 4307 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 12070 4307 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11988 4307 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11988 4307 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11906 4307 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11906 4307 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11824 4307 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11824 4307 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11742 4307 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11742 4307 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11660 4307 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11660 4307 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11578 4307 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11578 4307 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11496 4307 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11496 4307 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11414 4307 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11414 4307 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11332 4307 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11332 4307 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4243 11250 4307 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4243 11250 4307 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 12070 4226 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 12070 4226 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11988 4226 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11988 4226 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11906 4226 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11906 4226 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11824 4226 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11824 4226 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11742 4226 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11742 4226 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11660 4226 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11660 4226 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11578 4226 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11578 4226 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11496 4226 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11496 4226 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11414 4226 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11414 4226 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11332 4226 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11332 4226 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4162 11250 4226 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4162 11250 4226 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 12070 4145 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 12070 4145 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11988 4145 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11988 4145 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11906 4145 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11906 4145 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11824 4145 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11824 4145 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11742 4145 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11742 4145 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11660 4145 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11660 4145 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11578 4145 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11578 4145 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11496 4145 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11496 4145 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11414 4145 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11414 4145 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11332 4145 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11332 4145 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4081 11250 4145 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4081 11250 4145 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 12070 4064 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 12070 4064 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11988 4064 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11988 4064 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11906 4064 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11906 4064 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11824 4064 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11824 4064 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11742 4064 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11742 4064 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11660 4064 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11660 4064 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11578 4064 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11578 4064 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11496 4064 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11496 4064 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11414 4064 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11414 4064 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11332 4064 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11332 4064 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 4000 11250 4064 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 4000 11250 4064 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 12070 3983 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 12070 3983 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11988 3983 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11988 3983 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11906 3983 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11906 3983 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11824 3983 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11824 3983 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11742 3983 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11742 3983 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11660 3983 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11660 3983 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11578 3983 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11578 3983 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11496 3983 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11496 3983 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11414 3983 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11414 3983 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11332 3983 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11332 3983 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3919 11250 3983 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3919 11250 3983 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 12070 3902 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 12070 3902 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11988 3902 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11988 3902 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11906 3902 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11906 3902 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11824 3902 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11824 3902 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11742 3902 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11742 3902 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11660 3902 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11660 3902 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11578 3902 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11578 3902 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11496 3902 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11496 3902 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11414 3902 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11414 3902 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11332 3902 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11332 3902 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3838 11250 3902 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3838 11250 3902 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 12070 3821 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 12070 3821 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11988 3821 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11988 3821 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11906 3821 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11906 3821 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11824 3821 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11824 3821 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11742 3821 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11742 3821 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11660 3821 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11660 3821 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11578 3821 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11578 3821 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11496 3821 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11496 3821 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11414 3821 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11414 3821 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11332 3821 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11332 3821 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3757 11250 3821 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3757 11250 3821 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 12070 3740 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 12070 3740 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11988 3740 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11988 3740 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11906 3740 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11906 3740 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11824 3740 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11824 3740 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11742 3740 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11742 3740 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11660 3740 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11660 3740 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11578 3740 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11578 3740 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11496 3740 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11496 3740 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11414 3740 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11414 3740 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11332 3740 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11332 3740 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3676 11250 3740 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3676 11250 3740 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 12070 3659 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 12070 3659 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11988 3659 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11988 3659 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11906 3659 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11906 3659 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11824 3659 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11824 3659 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11742 3659 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11742 3659 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11660 3659 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11660 3659 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11578 3659 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11578 3659 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11496 3659 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11496 3659 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11414 3659 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11414 3659 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11332 3659 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11332 3659 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3595 11250 3659 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3595 11250 3659 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 12070 3578 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 12070 3578 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11988 3578 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11988 3578 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11906 3578 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11906 3578 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11824 3578 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11824 3578 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11742 3578 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11742 3578 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11660 3578 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11660 3578 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11578 3578 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11578 3578 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11496 3578 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11496 3578 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11414 3578 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11414 3578 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11332 3578 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11332 3578 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3514 11250 3578 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3514 11250 3578 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 12070 3497 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 12070 3497 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11988 3497 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11988 3497 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11906 3497 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11906 3497 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11824 3497 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11824 3497 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11742 3497 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11742 3497 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11660 3497 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11660 3497 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11578 3497 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11578 3497 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11496 3497 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11496 3497 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11414 3497 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11414 3497 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11332 3497 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11332 3497 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3433 11250 3497 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3433 11250 3497 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 12070 3416 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 12070 3416 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11988 3416 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11988 3416 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11906 3416 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11906 3416 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11824 3416 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11824 3416 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11742 3416 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11742 3416 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11660 3416 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11660 3416 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11578 3416 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11578 3416 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11496 3416 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11496 3416 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11414 3416 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11414 3416 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11332 3416 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11332 3416 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3352 11250 3416 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3352 11250 3416 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 12070 3335 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 12070 3335 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11988 3335 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11988 3335 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11906 3335 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11906 3335 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11824 3335 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11824 3335 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11742 3335 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11742 3335 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11660 3335 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11660 3335 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11578 3335 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11578 3335 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11496 3335 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11496 3335 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11414 3335 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11414 3335 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11332 3335 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11332 3335 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3271 11250 3335 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3271 11250 3335 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 12070 3254 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 12070 3254 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11988 3254 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11988 3254 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11906 3254 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11906 3254 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11824 3254 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11824 3254 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11742 3254 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11742 3254 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11660 3254 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11660 3254 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11578 3254 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11578 3254 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11496 3254 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11496 3254 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11414 3254 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11414 3254 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11332 3254 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11332 3254 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3190 11250 3254 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3190 11250 3254 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 12070 3173 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 12070 3173 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11988 3173 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11988 3173 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11906 3173 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11906 3173 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11824 3173 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11824 3173 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11742 3173 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11742 3173 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11660 3173 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11660 3173 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11578 3173 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11578 3173 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11496 3173 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11496 3173 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11414 3173 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11414 3173 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11332 3173 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11332 3173 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3109 11250 3173 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3109 11250 3173 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 12070 3092 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 12070 3092 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11988 3092 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11988 3092 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11906 3092 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11906 3092 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11824 3092 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11824 3092 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11742 3092 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11742 3092 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11660 3092 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11660 3092 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11578 3092 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11578 3092 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11496 3092 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11496 3092 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11414 3092 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11414 3092 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11332 3092 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11332 3092 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 3028 11250 3092 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 3028 11250 3092 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 12070 3011 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 12070 3011 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11988 3011 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11988 3011 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11906 3011 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11906 3011 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11824 3011 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11824 3011 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11742 3011 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11742 3011 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11660 3011 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11660 3011 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11578 3011 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11578 3011 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11496 3011 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11496 3011 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11414 3011 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11414 3011 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11332 3011 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11332 3011 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2947 11250 3011 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2947 11250 3011 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 12070 2930 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 12070 2930 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11988 2930 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11988 2930 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11906 2930 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11906 2930 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11824 2930 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11824 2930 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11742 2930 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11742 2930 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11660 2930 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11660 2930 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11578 2930 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11578 2930 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11496 2930 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11496 2930 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11414 2930 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11414 2930 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11332 2930 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11332 2930 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2866 11250 2930 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2866 11250 2930 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 12070 2849 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 12070 2849 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11988 2849 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11988 2849 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11906 2849 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11906 2849 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11824 2849 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11824 2849 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11742 2849 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11742 2849 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11660 2849 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11660 2849 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11578 2849 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11578 2849 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11496 2849 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11496 2849 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11414 2849 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11414 2849 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11332 2849 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11332 2849 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2785 11250 2849 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2785 11250 2849 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 12070 2768 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 12070 2768 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11988 2768 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11988 2768 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11906 2768 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11906 2768 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11824 2768 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11824 2768 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11742 2768 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11742 2768 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11660 2768 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11660 2768 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11578 2768 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11578 2768 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11496 2768 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11496 2768 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11414 2768 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11414 2768 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11332 2768 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11332 2768 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2704 11250 2768 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2704 11250 2768 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 12070 2687 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 12070 2687 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11988 2687 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11988 2687 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11906 2687 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11906 2687 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11824 2687 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11824 2687 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11742 2687 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11742 2687 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11660 2687 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11660 2687 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11578 2687 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11578 2687 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11496 2687 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11496 2687 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11414 2687 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11414 2687 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11332 2687 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11332 2687 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2623 11250 2687 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2623 11250 2687 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 12070 2606 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 12070 2606 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11988 2606 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11988 2606 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11906 2606 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11906 2606 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11824 2606 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11824 2606 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11742 2606 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11742 2606 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11660 2606 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11660 2606 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11578 2606 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11578 2606 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11496 2606 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11496 2606 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11414 2606 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11414 2606 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11332 2606 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11332 2606 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2542 11250 2606 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2542 11250 2606 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 12070 2525 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 12070 2525 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11988 2525 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11988 2525 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11906 2525 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11906 2525 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11824 2525 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11824 2525 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11742 2525 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11742 2525 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11660 2525 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11660 2525 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11578 2525 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11578 2525 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11496 2525 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11496 2525 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11414 2525 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11414 2525 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11332 2525 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11332 2525 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2461 11250 2525 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2461 11250 2525 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 12070 2444 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 12070 2444 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11988 2444 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11988 2444 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11906 2444 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11906 2444 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11824 2444 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11824 2444 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11742 2444 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11742 2444 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11660 2444 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11660 2444 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11578 2444 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11578 2444 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11496 2444 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11496 2444 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11414 2444 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11414 2444 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11332 2444 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11332 2444 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2380 11250 2444 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2380 11250 2444 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 12070 2363 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 12070 2363 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11988 2363 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11988 2363 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11906 2363 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11906 2363 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11824 2363 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11824 2363 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11742 2363 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11742 2363 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11660 2363 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11660 2363 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11578 2363 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11578 2363 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11496 2363 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11496 2363 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11414 2363 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11414 2363 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11332 2363 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11332 2363 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2299 11250 2363 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2299 11250 2363 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 12070 2282 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 12070 2282 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11988 2282 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11988 2282 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11906 2282 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11906 2282 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11824 2282 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11824 2282 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11742 2282 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11742 2282 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11660 2282 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11660 2282 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11578 2282 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11578 2282 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11496 2282 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11496 2282 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11414 2282 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11414 2282 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11332 2282 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11332 2282 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2218 11250 2282 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2218 11250 2282 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 12070 2201 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 12070 2201 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11988 2201 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11988 2201 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11906 2201 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11906 2201 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11824 2201 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11824 2201 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11742 2201 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11742 2201 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11660 2201 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11660 2201 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11578 2201 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11578 2201 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11496 2201 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11496 2201 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11414 2201 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11414 2201 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11332 2201 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11332 2201 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2137 11250 2201 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2137 11250 2201 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 12070 2120 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 12070 2120 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11988 2120 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11988 2120 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11906 2120 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11906 2120 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11824 2120 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11824 2120 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11742 2120 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11742 2120 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11660 2120 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11660 2120 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11578 2120 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11578 2120 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11496 2120 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11496 2120 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11414 2120 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11414 2120 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11332 2120 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11332 2120 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 2056 11250 2120 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 2056 11250 2120 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 12070 2039 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 12070 2039 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11988 2039 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11988 2039 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11906 2039 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11906 2039 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11824 2039 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11824 2039 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11742 2039 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11742 2039 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11660 2039 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11660 2039 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11578 2039 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11578 2039 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11496 2039 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11496 2039 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11414 2039 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11414 2039 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11332 2039 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11332 2039 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1975 11250 2039 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1975 11250 2039 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 12070 1958 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 12070 1958 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11988 1958 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11988 1958 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11906 1958 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11906 1958 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11824 1958 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11824 1958 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11742 1958 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11742 1958 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11660 1958 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11660 1958 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11578 1958 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11578 1958 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11496 1958 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11496 1958 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11414 1958 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11414 1958 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11332 1958 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11332 1958 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1894 11250 1958 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1894 11250 1958 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 12070 1877 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 12070 1877 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11988 1877 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11988 1877 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11906 1877 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11906 1877 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11824 1877 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11824 1877 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11742 1877 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11742 1877 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11660 1877 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11660 1877 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11578 1877 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11578 1877 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11496 1877 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11496 1877 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11414 1877 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11414 1877 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11332 1877 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11332 1877 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1813 11250 1877 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1813 11250 1877 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 12070 1796 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 12070 1796 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11988 1796 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11988 1796 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11906 1796 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11906 1796 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11824 1796 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11824 1796 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11742 1796 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11742 1796 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11660 1796 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11660 1796 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11578 1796 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11578 1796 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11496 1796 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11496 1796 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11414 1796 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11414 1796 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11332 1796 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11332 1796 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1732 11250 1796 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1732 11250 1796 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 12070 1715 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 12070 1715 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11988 1715 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11988 1715 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11906 1715 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11906 1715 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11824 1715 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11824 1715 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11742 1715 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11742 1715 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11660 1715 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11660 1715 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11578 1715 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11578 1715 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11496 1715 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11496 1715 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11414 1715 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11414 1715 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11332 1715 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11332 1715 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1651 11250 1715 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1651 11250 1715 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 12070 1634 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 12070 1634 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11988 1634 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11988 1634 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11906 1634 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11906 1634 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11824 1634 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11824 1634 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11742 1634 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11742 1634 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11660 1634 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11660 1634 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11578 1634 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11578 1634 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11496 1634 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11496 1634 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11414 1634 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11414 1634 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11332 1634 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11332 1634 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1570 11250 1634 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1570 11250 1634 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 12070 1553 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 12070 1553 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11988 1553 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11988 1553 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11906 1553 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11906 1553 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11824 1553 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11824 1553 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11742 1553 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11742 1553 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11660 1553 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11660 1553 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11578 1553 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11578 1553 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11496 1553 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11496 1553 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11414 1553 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11414 1553 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11332 1553 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11332 1553 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1489 11250 1553 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1489 11250 1553 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 12070 1472 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 12070 1472 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11988 1472 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11988 1472 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11906 1472 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11906 1472 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11824 1472 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11824 1472 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11742 1472 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11742 1472 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11660 1472 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11660 1472 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11578 1472 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11578 1472 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11496 1472 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11496 1472 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11414 1472 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11414 1472 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11332 1472 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11332 1472 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1408 11250 1472 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1408 11250 1472 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 12070 1391 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 12070 1391 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11988 1391 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11988 1391 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11906 1391 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11906 1391 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11824 1391 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11824 1391 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11742 1391 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11742 1391 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11660 1391 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11660 1391 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11578 1391 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11578 1391 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11496 1391 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11496 1391 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11414 1391 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11414 1391 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11332 1391 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11332 1391 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1327 11250 1391 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1327 11250 1391 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 12070 1310 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 12070 1310 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11988 1310 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11988 1310 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11906 1310 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11906 1310 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11824 1310 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11824 1310 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11742 1310 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11742 1310 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11660 1310 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11660 1310 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11578 1310 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11578 1310 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11496 1310 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11496 1310 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11414 1310 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11414 1310 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11332 1310 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11332 1310 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1246 11250 1310 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1246 11250 1310 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 12070 1229 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 12070 1229 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11988 1229 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11988 1229 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11906 1229 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11906 1229 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11824 1229 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11824 1229 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11742 1229 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11742 1229 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11660 1229 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11660 1229 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11578 1229 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11578 1229 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11496 1229 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11496 1229 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11414 1229 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11414 1229 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11332 1229 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11332 1229 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1165 11250 1229 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1165 11250 1229 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 12070 1148 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 12070 1148 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11988 1148 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11988 1148 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11906 1148 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11906 1148 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11824 1148 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11824 1148 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11742 1148 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11742 1148 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11660 1148 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11660 1148 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11578 1148 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11578 1148 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11496 1148 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11496 1148 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11414 1148 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11414 1148 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11332 1148 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11332 1148 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1084 11250 1148 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1084 11250 1148 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 12070 1067 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 12070 1067 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11988 1067 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11988 1067 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11906 1067 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11906 1067 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11824 1067 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11824 1067 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11742 1067 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11742 1067 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11660 1067 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11660 1067 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11578 1067 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11578 1067 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11496 1067 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11496 1067 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11414 1067 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11414 1067 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11332 1067 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11332 1067 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 1003 11250 1067 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 1003 11250 1067 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 12070 986 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 12070 986 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11988 986 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11988 986 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11906 986 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11906 986 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11824 986 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11824 986 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11742 986 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11742 986 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11660 986 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11660 986 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11578 986 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11578 986 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11496 986 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11496 986 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11414 986 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11414 986 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11332 986 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11332 986 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 922 11250 986 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 922 11250 986 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 12070 905 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 12070 905 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11988 905 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11988 905 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11906 905 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11906 905 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11824 905 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11824 905 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11742 905 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11742 905 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11660 905 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11660 905 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11578 905 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11578 905 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11496 905 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11496 905 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11414 905 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11414 905 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11332 905 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11332 905 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 841 11250 905 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 841 11250 905 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 12070 824 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 12070 824 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11988 824 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11988 824 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11906 824 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11906 824 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11824 824 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11824 824 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11742 824 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11742 824 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11660 824 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11660 824 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11578 824 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11578 824 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11496 824 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11496 824 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11414 824 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11414 824 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11332 824 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11332 824 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 760 11250 824 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 760 11250 824 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 12070 743 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 12070 743 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11988 743 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11988 743 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11906 743 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11906 743 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11824 743 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11824 743 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11742 743 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11742 743 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11660 743 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11660 743 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11578 743 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11578 743 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11496 743 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11496 743 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11414 743 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11414 743 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11332 743 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11332 743 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 679 11250 743 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 679 11250 743 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 12070 662 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 12070 662 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11988 662 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11988 662 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11906 662 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11906 662 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11824 662 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11824 662 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11742 662 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11742 662 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11660 662 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11660 662 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11578 662 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11578 662 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11496 662 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11496 662 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11414 662 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11414 662 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11332 662 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11332 662 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 598 11250 662 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 598 11250 662 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 12070 580 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 12070 580 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11988 580 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11988 580 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11906 580 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11906 580 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11824 580 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11824 580 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11742 580 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11742 580 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11660 580 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11660 580 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11578 580 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11578 580 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11496 580 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11496 580 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11414 580 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11414 580 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11332 580 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11332 580 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 516 11250 580 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 516 11250 580 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 12070 498 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 12070 498 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11988 498 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11988 498 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11906 498 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11906 498 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11824 498 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11824 498 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11742 498 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11742 498 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11660 498 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11660 498 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11578 498 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11578 498 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11496 498 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11496 498 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11414 498 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11414 498 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11332 498 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11332 498 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 434 11250 498 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 434 11250 498 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 12070 416 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 12070 416 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11988 416 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11988 416 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11906 416 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11906 416 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11824 416 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11824 416 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11742 416 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11742 416 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11660 416 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11660 416 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11578 416 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11578 416 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11496 416 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11496 416 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11414 416 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11414 416 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11332 416 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11332 416 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 352 11250 416 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 352 11250 416 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 12070 334 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 12070 334 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11988 334 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11988 334 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11906 334 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11906 334 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11824 334 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11824 334 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11742 334 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11742 334 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11660 334 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11660 334 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11578 334 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11578 334 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11496 334 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11496 334 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11414 334 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11414 334 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11332 334 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11332 334 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 270 11250 334 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 270 11250 334 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 12070 252 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11988 252 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11906 252 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11824 252 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11742 252 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11660 252 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11578 252 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11496 252 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11414 252 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11332 252 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 188 11250 252 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 12070 170 12134 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11988 170 12052 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11906 170 11970 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11824 170 11888 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11742 170 11806 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11660 170 11724 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11578 170 11642 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11496 170 11560 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11414 170 11478 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11332 170 11396 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal3 s 106 11250 170 11314 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 57 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 58 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 59 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 60 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 60 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 60 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 60 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 24961536
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 24549616
<< end >>
