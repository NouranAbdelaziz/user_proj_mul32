/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hvl/cdl/sky130_fd_sc_hvl.cdl