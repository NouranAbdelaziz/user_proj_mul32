/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/klayout/pymacros/cells/fixed_devices/VPP/sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4.cdl