magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< pwell >>
rect 10 66 1014 1536
<< mvnmos >>
rect 228 92 328 1510
rect 384 92 484 1510
rect 540 92 640 1510
rect 696 92 796 1510
<< mvndiff >>
rect 172 1498 228 1510
rect 172 1464 183 1498
rect 217 1464 228 1498
rect 172 1430 228 1464
rect 172 1396 183 1430
rect 217 1396 228 1430
rect 172 1362 228 1396
rect 172 1328 183 1362
rect 217 1328 228 1362
rect 172 1294 228 1328
rect 172 1260 183 1294
rect 217 1260 228 1294
rect 172 1226 228 1260
rect 172 1192 183 1226
rect 217 1192 228 1226
rect 172 1158 228 1192
rect 172 1124 183 1158
rect 217 1124 228 1158
rect 172 1090 228 1124
rect 172 1056 183 1090
rect 217 1056 228 1090
rect 172 1022 228 1056
rect 172 988 183 1022
rect 217 988 228 1022
rect 172 954 228 988
rect 172 920 183 954
rect 217 920 228 954
rect 172 886 228 920
rect 172 852 183 886
rect 217 852 228 886
rect 172 818 228 852
rect 172 784 183 818
rect 217 784 228 818
rect 172 750 228 784
rect 172 716 183 750
rect 217 716 228 750
rect 172 682 228 716
rect 172 648 183 682
rect 217 648 228 682
rect 172 614 228 648
rect 172 580 183 614
rect 217 580 228 614
rect 172 546 228 580
rect 172 512 183 546
rect 217 512 228 546
rect 172 478 228 512
rect 172 444 183 478
rect 217 444 228 478
rect 172 410 228 444
rect 172 376 183 410
rect 217 376 228 410
rect 172 342 228 376
rect 172 308 183 342
rect 217 308 228 342
rect 172 274 228 308
rect 172 240 183 274
rect 217 240 228 274
rect 172 206 228 240
rect 172 172 183 206
rect 217 172 228 206
rect 172 138 228 172
rect 172 104 183 138
rect 217 104 228 138
rect 172 92 228 104
rect 328 1498 384 1510
rect 328 1464 339 1498
rect 373 1464 384 1498
rect 328 1430 384 1464
rect 328 1396 339 1430
rect 373 1396 384 1430
rect 328 1362 384 1396
rect 328 1328 339 1362
rect 373 1328 384 1362
rect 328 1294 384 1328
rect 328 1260 339 1294
rect 373 1260 384 1294
rect 328 1226 384 1260
rect 328 1192 339 1226
rect 373 1192 384 1226
rect 328 1158 384 1192
rect 328 1124 339 1158
rect 373 1124 384 1158
rect 328 1090 384 1124
rect 328 1056 339 1090
rect 373 1056 384 1090
rect 328 1022 384 1056
rect 328 988 339 1022
rect 373 988 384 1022
rect 328 954 384 988
rect 328 920 339 954
rect 373 920 384 954
rect 328 886 384 920
rect 328 852 339 886
rect 373 852 384 886
rect 328 818 384 852
rect 328 784 339 818
rect 373 784 384 818
rect 328 750 384 784
rect 328 716 339 750
rect 373 716 384 750
rect 328 682 384 716
rect 328 648 339 682
rect 373 648 384 682
rect 328 614 384 648
rect 328 580 339 614
rect 373 580 384 614
rect 328 546 384 580
rect 328 512 339 546
rect 373 512 384 546
rect 328 478 384 512
rect 328 444 339 478
rect 373 444 384 478
rect 328 410 384 444
rect 328 376 339 410
rect 373 376 384 410
rect 328 342 384 376
rect 328 308 339 342
rect 373 308 384 342
rect 328 274 384 308
rect 328 240 339 274
rect 373 240 384 274
rect 328 206 384 240
rect 328 172 339 206
rect 373 172 384 206
rect 328 138 384 172
rect 328 104 339 138
rect 373 104 384 138
rect 328 92 384 104
rect 484 1498 540 1510
rect 484 1464 495 1498
rect 529 1464 540 1498
rect 484 1430 540 1464
rect 484 1396 495 1430
rect 529 1396 540 1430
rect 484 1362 540 1396
rect 484 1328 495 1362
rect 529 1328 540 1362
rect 484 1294 540 1328
rect 484 1260 495 1294
rect 529 1260 540 1294
rect 484 1226 540 1260
rect 484 1192 495 1226
rect 529 1192 540 1226
rect 484 1158 540 1192
rect 484 1124 495 1158
rect 529 1124 540 1158
rect 484 1090 540 1124
rect 484 1056 495 1090
rect 529 1056 540 1090
rect 484 1022 540 1056
rect 484 988 495 1022
rect 529 988 540 1022
rect 484 954 540 988
rect 484 920 495 954
rect 529 920 540 954
rect 484 886 540 920
rect 484 852 495 886
rect 529 852 540 886
rect 484 818 540 852
rect 484 784 495 818
rect 529 784 540 818
rect 484 750 540 784
rect 484 716 495 750
rect 529 716 540 750
rect 484 682 540 716
rect 484 648 495 682
rect 529 648 540 682
rect 484 614 540 648
rect 484 580 495 614
rect 529 580 540 614
rect 484 546 540 580
rect 484 512 495 546
rect 529 512 540 546
rect 484 478 540 512
rect 484 444 495 478
rect 529 444 540 478
rect 484 410 540 444
rect 484 376 495 410
rect 529 376 540 410
rect 484 342 540 376
rect 484 308 495 342
rect 529 308 540 342
rect 484 274 540 308
rect 484 240 495 274
rect 529 240 540 274
rect 484 206 540 240
rect 484 172 495 206
rect 529 172 540 206
rect 484 138 540 172
rect 484 104 495 138
rect 529 104 540 138
rect 484 92 540 104
rect 640 1498 696 1510
rect 640 1464 651 1498
rect 685 1464 696 1498
rect 640 1430 696 1464
rect 640 1396 651 1430
rect 685 1396 696 1430
rect 640 1362 696 1396
rect 640 1328 651 1362
rect 685 1328 696 1362
rect 640 1294 696 1328
rect 640 1260 651 1294
rect 685 1260 696 1294
rect 640 1226 696 1260
rect 640 1192 651 1226
rect 685 1192 696 1226
rect 640 1158 696 1192
rect 640 1124 651 1158
rect 685 1124 696 1158
rect 640 1090 696 1124
rect 640 1056 651 1090
rect 685 1056 696 1090
rect 640 1022 696 1056
rect 640 988 651 1022
rect 685 988 696 1022
rect 640 954 696 988
rect 640 920 651 954
rect 685 920 696 954
rect 640 886 696 920
rect 640 852 651 886
rect 685 852 696 886
rect 640 818 696 852
rect 640 784 651 818
rect 685 784 696 818
rect 640 750 696 784
rect 640 716 651 750
rect 685 716 696 750
rect 640 682 696 716
rect 640 648 651 682
rect 685 648 696 682
rect 640 614 696 648
rect 640 580 651 614
rect 685 580 696 614
rect 640 546 696 580
rect 640 512 651 546
rect 685 512 696 546
rect 640 478 696 512
rect 640 444 651 478
rect 685 444 696 478
rect 640 410 696 444
rect 640 376 651 410
rect 685 376 696 410
rect 640 342 696 376
rect 640 308 651 342
rect 685 308 696 342
rect 640 274 696 308
rect 640 240 651 274
rect 685 240 696 274
rect 640 206 696 240
rect 640 172 651 206
rect 685 172 696 206
rect 640 138 696 172
rect 640 104 651 138
rect 685 104 696 138
rect 640 92 696 104
rect 796 1498 852 1510
rect 796 1464 807 1498
rect 841 1464 852 1498
rect 796 1430 852 1464
rect 796 1396 807 1430
rect 841 1396 852 1430
rect 796 1362 852 1396
rect 796 1328 807 1362
rect 841 1328 852 1362
rect 796 1294 852 1328
rect 796 1260 807 1294
rect 841 1260 852 1294
rect 796 1226 852 1260
rect 796 1192 807 1226
rect 841 1192 852 1226
rect 796 1158 852 1192
rect 796 1124 807 1158
rect 841 1124 852 1158
rect 796 1090 852 1124
rect 796 1056 807 1090
rect 841 1056 852 1090
rect 796 1022 852 1056
rect 796 988 807 1022
rect 841 988 852 1022
rect 796 954 852 988
rect 796 920 807 954
rect 841 920 852 954
rect 796 886 852 920
rect 796 852 807 886
rect 841 852 852 886
rect 796 818 852 852
rect 796 784 807 818
rect 841 784 852 818
rect 796 750 852 784
rect 796 716 807 750
rect 841 716 852 750
rect 796 682 852 716
rect 796 648 807 682
rect 841 648 852 682
rect 796 614 852 648
rect 796 580 807 614
rect 841 580 852 614
rect 796 546 852 580
rect 796 512 807 546
rect 841 512 852 546
rect 796 478 852 512
rect 796 444 807 478
rect 841 444 852 478
rect 796 410 852 444
rect 796 376 807 410
rect 841 376 852 410
rect 796 342 852 376
rect 796 308 807 342
rect 841 308 852 342
rect 796 274 852 308
rect 796 240 807 274
rect 841 240 852 274
rect 796 206 852 240
rect 796 172 807 206
rect 841 172 852 206
rect 796 138 852 172
rect 796 104 807 138
rect 841 104 852 138
rect 796 92 852 104
<< mvndiffc >>
rect 183 1464 217 1498
rect 183 1396 217 1430
rect 183 1328 217 1362
rect 183 1260 217 1294
rect 183 1192 217 1226
rect 183 1124 217 1158
rect 183 1056 217 1090
rect 183 988 217 1022
rect 183 920 217 954
rect 183 852 217 886
rect 183 784 217 818
rect 183 716 217 750
rect 183 648 217 682
rect 183 580 217 614
rect 183 512 217 546
rect 183 444 217 478
rect 183 376 217 410
rect 183 308 217 342
rect 183 240 217 274
rect 183 172 217 206
rect 183 104 217 138
rect 339 1464 373 1498
rect 339 1396 373 1430
rect 339 1328 373 1362
rect 339 1260 373 1294
rect 339 1192 373 1226
rect 339 1124 373 1158
rect 339 1056 373 1090
rect 339 988 373 1022
rect 339 920 373 954
rect 339 852 373 886
rect 339 784 373 818
rect 339 716 373 750
rect 339 648 373 682
rect 339 580 373 614
rect 339 512 373 546
rect 339 444 373 478
rect 339 376 373 410
rect 339 308 373 342
rect 339 240 373 274
rect 339 172 373 206
rect 339 104 373 138
rect 495 1464 529 1498
rect 495 1396 529 1430
rect 495 1328 529 1362
rect 495 1260 529 1294
rect 495 1192 529 1226
rect 495 1124 529 1158
rect 495 1056 529 1090
rect 495 988 529 1022
rect 495 920 529 954
rect 495 852 529 886
rect 495 784 529 818
rect 495 716 529 750
rect 495 648 529 682
rect 495 580 529 614
rect 495 512 529 546
rect 495 444 529 478
rect 495 376 529 410
rect 495 308 529 342
rect 495 240 529 274
rect 495 172 529 206
rect 495 104 529 138
rect 651 1464 685 1498
rect 651 1396 685 1430
rect 651 1328 685 1362
rect 651 1260 685 1294
rect 651 1192 685 1226
rect 651 1124 685 1158
rect 651 1056 685 1090
rect 651 988 685 1022
rect 651 920 685 954
rect 651 852 685 886
rect 651 784 685 818
rect 651 716 685 750
rect 651 648 685 682
rect 651 580 685 614
rect 651 512 685 546
rect 651 444 685 478
rect 651 376 685 410
rect 651 308 685 342
rect 651 240 685 274
rect 651 172 685 206
rect 651 104 685 138
rect 807 1464 841 1498
rect 807 1396 841 1430
rect 807 1328 841 1362
rect 807 1260 841 1294
rect 807 1192 841 1226
rect 807 1124 841 1158
rect 807 1056 841 1090
rect 807 988 841 1022
rect 807 920 841 954
rect 807 852 841 886
rect 807 784 841 818
rect 807 716 841 750
rect 807 648 841 682
rect 807 580 841 614
rect 807 512 841 546
rect 807 444 841 478
rect 807 376 841 410
rect 807 308 841 342
rect 807 240 841 274
rect 807 172 841 206
rect 807 104 841 138
<< mvpsubdiff >>
rect 36 1464 94 1510
rect 36 1430 48 1464
rect 82 1430 94 1464
rect 36 1396 94 1430
rect 36 1362 48 1396
rect 82 1362 94 1396
rect 36 1328 94 1362
rect 36 1294 48 1328
rect 82 1294 94 1328
rect 36 1260 94 1294
rect 36 1226 48 1260
rect 82 1226 94 1260
rect 36 1192 94 1226
rect 36 1158 48 1192
rect 82 1158 94 1192
rect 36 1124 94 1158
rect 36 1090 48 1124
rect 82 1090 94 1124
rect 36 1056 94 1090
rect 36 1022 48 1056
rect 82 1022 94 1056
rect 36 988 94 1022
rect 36 954 48 988
rect 82 954 94 988
rect 36 920 94 954
rect 36 886 48 920
rect 82 886 94 920
rect 36 852 94 886
rect 36 818 48 852
rect 82 818 94 852
rect 36 784 94 818
rect 36 750 48 784
rect 82 750 94 784
rect 36 716 94 750
rect 36 682 48 716
rect 82 682 94 716
rect 36 648 94 682
rect 36 614 48 648
rect 82 614 94 648
rect 36 580 94 614
rect 36 546 48 580
rect 82 546 94 580
rect 36 512 94 546
rect 36 478 48 512
rect 82 478 94 512
rect 36 444 94 478
rect 36 410 48 444
rect 82 410 94 444
rect 36 376 94 410
rect 36 342 48 376
rect 82 342 94 376
rect 36 308 94 342
rect 36 274 48 308
rect 82 274 94 308
rect 36 240 94 274
rect 36 206 48 240
rect 82 206 94 240
rect 36 172 94 206
rect 36 138 48 172
rect 82 138 94 172
rect 36 92 94 138
rect 930 1464 988 1510
rect 930 1430 942 1464
rect 976 1430 988 1464
rect 930 1396 988 1430
rect 930 1362 942 1396
rect 976 1362 988 1396
rect 930 1328 988 1362
rect 930 1294 942 1328
rect 976 1294 988 1328
rect 930 1260 988 1294
rect 930 1226 942 1260
rect 976 1226 988 1260
rect 930 1192 988 1226
rect 930 1158 942 1192
rect 976 1158 988 1192
rect 930 1124 988 1158
rect 930 1090 942 1124
rect 976 1090 988 1124
rect 930 1056 988 1090
rect 930 1022 942 1056
rect 976 1022 988 1056
rect 930 988 988 1022
rect 930 954 942 988
rect 976 954 988 988
rect 930 920 988 954
rect 930 886 942 920
rect 976 886 988 920
rect 930 852 988 886
rect 930 818 942 852
rect 976 818 988 852
rect 930 784 988 818
rect 930 750 942 784
rect 976 750 988 784
rect 930 716 988 750
rect 930 682 942 716
rect 976 682 988 716
rect 930 648 988 682
rect 930 614 942 648
rect 976 614 988 648
rect 930 580 988 614
rect 930 546 942 580
rect 976 546 988 580
rect 930 512 988 546
rect 930 478 942 512
rect 976 478 988 512
rect 930 444 988 478
rect 930 410 942 444
rect 976 410 988 444
rect 930 376 988 410
rect 930 342 942 376
rect 976 342 988 376
rect 930 308 988 342
rect 930 274 942 308
rect 976 274 988 308
rect 930 240 988 274
rect 930 206 942 240
rect 976 206 988 240
rect 930 172 988 206
rect 930 138 942 172
rect 976 138 988 172
rect 930 92 988 138
<< mvpsubdiffcont >>
rect 48 1430 82 1464
rect 48 1362 82 1396
rect 48 1294 82 1328
rect 48 1226 82 1260
rect 48 1158 82 1192
rect 48 1090 82 1124
rect 48 1022 82 1056
rect 48 954 82 988
rect 48 886 82 920
rect 48 818 82 852
rect 48 750 82 784
rect 48 682 82 716
rect 48 614 82 648
rect 48 546 82 580
rect 48 478 82 512
rect 48 410 82 444
rect 48 342 82 376
rect 48 274 82 308
rect 48 206 82 240
rect 48 138 82 172
rect 942 1430 976 1464
rect 942 1362 976 1396
rect 942 1294 976 1328
rect 942 1226 976 1260
rect 942 1158 976 1192
rect 942 1090 976 1124
rect 942 1022 976 1056
rect 942 954 976 988
rect 942 886 976 920
rect 942 818 976 852
rect 942 750 976 784
rect 942 682 976 716
rect 942 614 976 648
rect 942 546 976 580
rect 942 478 976 512
rect 942 410 976 444
rect 942 342 976 376
rect 942 274 976 308
rect 942 206 976 240
rect 942 138 976 172
<< poly >>
rect 207 1582 817 1602
rect 207 1548 223 1582
rect 257 1548 291 1582
rect 325 1548 359 1582
rect 393 1548 427 1582
rect 461 1548 495 1582
rect 529 1548 563 1582
rect 597 1548 631 1582
rect 665 1548 699 1582
rect 733 1548 767 1582
rect 801 1548 817 1582
rect 207 1532 817 1548
rect 228 1510 328 1532
rect 384 1510 484 1532
rect 540 1510 640 1532
rect 696 1510 796 1532
rect 228 70 328 92
rect 384 70 484 92
rect 540 70 640 92
rect 696 70 796 92
rect 207 54 817 70
rect 207 20 223 54
rect 257 20 291 54
rect 325 20 359 54
rect 393 20 427 54
rect 461 20 495 54
rect 529 20 563 54
rect 597 20 631 54
rect 665 20 699 54
rect 733 20 767 54
rect 801 20 817 54
rect 207 0 817 20
<< polycont >>
rect 223 1548 257 1582
rect 291 1548 325 1582
rect 359 1548 393 1582
rect 427 1548 461 1582
rect 495 1548 529 1582
rect 563 1548 597 1582
rect 631 1548 665 1582
rect 699 1548 733 1582
rect 767 1548 801 1582
rect 223 20 257 54
rect 291 20 325 54
rect 359 20 393 54
rect 427 20 461 54
rect 495 20 529 54
rect 563 20 597 54
rect 631 20 665 54
rect 699 20 733 54
rect 767 20 801 54
<< locali >>
rect 207 1548 223 1582
rect 277 1548 291 1582
rect 349 1548 359 1582
rect 421 1548 427 1582
rect 493 1548 495 1582
rect 529 1548 531 1582
rect 597 1548 603 1582
rect 665 1548 675 1582
rect 733 1548 747 1582
rect 801 1548 817 1582
rect 48 1466 82 1514
rect 48 1396 82 1430
rect 48 1328 82 1360
rect 48 1260 82 1288
rect 48 1192 82 1216
rect 48 1124 82 1144
rect 48 1056 82 1072
rect 48 988 82 1000
rect 48 920 82 928
rect 48 852 82 856
rect 48 746 82 750
rect 48 674 82 682
rect 48 602 82 614
rect 48 530 82 546
rect 48 458 82 478
rect 48 386 82 410
rect 48 314 82 342
rect 48 242 82 274
rect 48 172 82 206
rect 48 88 82 136
rect 183 1498 217 1514
rect 183 1430 217 1432
rect 183 1394 217 1396
rect 183 1322 217 1328
rect 183 1250 217 1260
rect 183 1178 217 1192
rect 183 1106 217 1124
rect 183 1034 217 1056
rect 183 962 217 988
rect 183 890 217 920
rect 183 818 217 852
rect 183 750 217 784
rect 183 682 217 712
rect 183 614 217 640
rect 183 546 217 568
rect 183 478 217 496
rect 183 410 217 424
rect 183 342 217 352
rect 183 274 217 280
rect 183 206 217 208
rect 183 170 217 172
rect 183 88 217 104
rect 339 1498 373 1514
rect 339 1430 373 1432
rect 339 1394 373 1396
rect 339 1322 373 1328
rect 339 1250 373 1260
rect 339 1178 373 1192
rect 339 1106 373 1124
rect 339 1034 373 1056
rect 339 962 373 988
rect 339 890 373 920
rect 339 818 373 852
rect 339 750 373 784
rect 339 682 373 712
rect 339 614 373 640
rect 339 546 373 568
rect 339 478 373 496
rect 339 410 373 424
rect 339 342 373 352
rect 339 274 373 280
rect 339 206 373 208
rect 339 170 373 172
rect 339 88 373 104
rect 495 1498 529 1514
rect 495 1430 529 1432
rect 495 1394 529 1396
rect 495 1322 529 1328
rect 495 1250 529 1260
rect 495 1178 529 1192
rect 495 1106 529 1124
rect 495 1034 529 1056
rect 495 962 529 988
rect 495 890 529 920
rect 495 818 529 852
rect 495 750 529 784
rect 495 682 529 712
rect 495 614 529 640
rect 495 546 529 568
rect 495 478 529 496
rect 495 410 529 424
rect 495 342 529 352
rect 495 274 529 280
rect 495 206 529 208
rect 495 170 529 172
rect 495 88 529 104
rect 651 1498 685 1514
rect 651 1430 685 1432
rect 651 1394 685 1396
rect 651 1322 685 1328
rect 651 1250 685 1260
rect 651 1178 685 1192
rect 651 1106 685 1124
rect 651 1034 685 1056
rect 651 962 685 988
rect 651 890 685 920
rect 651 818 685 852
rect 651 750 685 784
rect 651 682 685 712
rect 651 614 685 640
rect 651 546 685 568
rect 651 478 685 496
rect 651 410 685 424
rect 651 342 685 352
rect 651 274 685 280
rect 651 206 685 208
rect 651 170 685 172
rect 651 88 685 104
rect 807 1498 841 1514
rect 807 1430 841 1432
rect 807 1394 841 1396
rect 807 1322 841 1328
rect 807 1250 841 1260
rect 807 1178 841 1192
rect 807 1106 841 1124
rect 807 1034 841 1056
rect 807 962 841 988
rect 807 890 841 920
rect 807 818 841 852
rect 807 750 841 784
rect 807 682 841 712
rect 807 614 841 640
rect 807 546 841 568
rect 807 478 841 496
rect 807 410 841 424
rect 807 342 841 352
rect 807 274 841 280
rect 807 206 841 208
rect 807 170 841 172
rect 942 1466 976 1480
rect 942 1396 976 1430
rect 942 1328 976 1360
rect 942 1260 976 1288
rect 942 1192 976 1216
rect 942 1124 976 1144
rect 942 1056 976 1072
rect 942 988 976 1000
rect 942 920 976 928
rect 942 852 976 856
rect 942 746 976 750
rect 942 674 976 682
rect 942 602 976 614
rect 942 530 976 546
rect 942 458 976 478
rect 942 386 976 410
rect 942 314 976 342
rect 942 242 976 274
rect 942 172 976 206
rect 942 122 976 136
rect 807 88 841 104
rect 207 20 223 54
rect 277 20 291 54
rect 349 20 359 54
rect 421 20 427 54
rect 493 20 495 54
rect 529 20 531 54
rect 597 20 603 54
rect 665 20 675 54
rect 733 20 747 54
rect 801 20 817 54
<< viali >>
rect 243 1548 257 1582
rect 257 1548 277 1582
rect 315 1548 325 1582
rect 325 1548 349 1582
rect 387 1548 393 1582
rect 393 1548 421 1582
rect 459 1548 461 1582
rect 461 1548 493 1582
rect 531 1548 563 1582
rect 563 1548 565 1582
rect 603 1548 631 1582
rect 631 1548 637 1582
rect 675 1548 699 1582
rect 699 1548 709 1582
rect 747 1548 767 1582
rect 767 1548 781 1582
rect 48 1464 82 1466
rect 48 1432 82 1464
rect 48 1362 82 1394
rect 48 1360 82 1362
rect 48 1294 82 1322
rect 48 1288 82 1294
rect 48 1226 82 1250
rect 48 1216 82 1226
rect 48 1158 82 1178
rect 48 1144 82 1158
rect 48 1090 82 1106
rect 48 1072 82 1090
rect 48 1022 82 1034
rect 48 1000 82 1022
rect 48 954 82 962
rect 48 928 82 954
rect 48 886 82 890
rect 48 856 82 886
rect 48 784 82 818
rect 48 716 82 746
rect 48 712 82 716
rect 48 648 82 674
rect 48 640 82 648
rect 48 580 82 602
rect 48 568 82 580
rect 48 512 82 530
rect 48 496 82 512
rect 48 444 82 458
rect 48 424 82 444
rect 48 376 82 386
rect 48 352 82 376
rect 48 308 82 314
rect 48 280 82 308
rect 48 240 82 242
rect 48 208 82 240
rect 48 138 82 170
rect 48 136 82 138
rect 183 1464 217 1466
rect 183 1432 217 1464
rect 183 1362 217 1394
rect 183 1360 217 1362
rect 183 1294 217 1322
rect 183 1288 217 1294
rect 183 1226 217 1250
rect 183 1216 217 1226
rect 183 1158 217 1178
rect 183 1144 217 1158
rect 183 1090 217 1106
rect 183 1072 217 1090
rect 183 1022 217 1034
rect 183 1000 217 1022
rect 183 954 217 962
rect 183 928 217 954
rect 183 886 217 890
rect 183 856 217 886
rect 183 784 217 818
rect 183 716 217 746
rect 183 712 217 716
rect 183 648 217 674
rect 183 640 217 648
rect 183 580 217 602
rect 183 568 217 580
rect 183 512 217 530
rect 183 496 217 512
rect 183 444 217 458
rect 183 424 217 444
rect 183 376 217 386
rect 183 352 217 376
rect 183 308 217 314
rect 183 280 217 308
rect 183 240 217 242
rect 183 208 217 240
rect 183 138 217 170
rect 183 136 217 138
rect 339 1464 373 1466
rect 339 1432 373 1464
rect 339 1362 373 1394
rect 339 1360 373 1362
rect 339 1294 373 1322
rect 339 1288 373 1294
rect 339 1226 373 1250
rect 339 1216 373 1226
rect 339 1158 373 1178
rect 339 1144 373 1158
rect 339 1090 373 1106
rect 339 1072 373 1090
rect 339 1022 373 1034
rect 339 1000 373 1022
rect 339 954 373 962
rect 339 928 373 954
rect 339 886 373 890
rect 339 856 373 886
rect 339 784 373 818
rect 339 716 373 746
rect 339 712 373 716
rect 339 648 373 674
rect 339 640 373 648
rect 339 580 373 602
rect 339 568 373 580
rect 339 512 373 530
rect 339 496 373 512
rect 339 444 373 458
rect 339 424 373 444
rect 339 376 373 386
rect 339 352 373 376
rect 339 308 373 314
rect 339 280 373 308
rect 339 240 373 242
rect 339 208 373 240
rect 339 138 373 170
rect 339 136 373 138
rect 495 1464 529 1466
rect 495 1432 529 1464
rect 495 1362 529 1394
rect 495 1360 529 1362
rect 495 1294 529 1322
rect 495 1288 529 1294
rect 495 1226 529 1250
rect 495 1216 529 1226
rect 495 1158 529 1178
rect 495 1144 529 1158
rect 495 1090 529 1106
rect 495 1072 529 1090
rect 495 1022 529 1034
rect 495 1000 529 1022
rect 495 954 529 962
rect 495 928 529 954
rect 495 886 529 890
rect 495 856 529 886
rect 495 784 529 818
rect 495 716 529 746
rect 495 712 529 716
rect 495 648 529 674
rect 495 640 529 648
rect 495 580 529 602
rect 495 568 529 580
rect 495 512 529 530
rect 495 496 529 512
rect 495 444 529 458
rect 495 424 529 444
rect 495 376 529 386
rect 495 352 529 376
rect 495 308 529 314
rect 495 280 529 308
rect 495 240 529 242
rect 495 208 529 240
rect 495 138 529 170
rect 495 136 529 138
rect 651 1464 685 1466
rect 651 1432 685 1464
rect 651 1362 685 1394
rect 651 1360 685 1362
rect 651 1294 685 1322
rect 651 1288 685 1294
rect 651 1226 685 1250
rect 651 1216 685 1226
rect 651 1158 685 1178
rect 651 1144 685 1158
rect 651 1090 685 1106
rect 651 1072 685 1090
rect 651 1022 685 1034
rect 651 1000 685 1022
rect 651 954 685 962
rect 651 928 685 954
rect 651 886 685 890
rect 651 856 685 886
rect 651 784 685 818
rect 651 716 685 746
rect 651 712 685 716
rect 651 648 685 674
rect 651 640 685 648
rect 651 580 685 602
rect 651 568 685 580
rect 651 512 685 530
rect 651 496 685 512
rect 651 444 685 458
rect 651 424 685 444
rect 651 376 685 386
rect 651 352 685 376
rect 651 308 685 314
rect 651 280 685 308
rect 651 240 685 242
rect 651 208 685 240
rect 651 138 685 170
rect 651 136 685 138
rect 807 1464 841 1466
rect 807 1432 841 1464
rect 807 1362 841 1394
rect 807 1360 841 1362
rect 807 1294 841 1322
rect 807 1288 841 1294
rect 807 1226 841 1250
rect 807 1216 841 1226
rect 807 1158 841 1178
rect 807 1144 841 1158
rect 807 1090 841 1106
rect 807 1072 841 1090
rect 807 1022 841 1034
rect 807 1000 841 1022
rect 807 954 841 962
rect 807 928 841 954
rect 807 886 841 890
rect 807 856 841 886
rect 807 784 841 818
rect 807 716 841 746
rect 807 712 841 716
rect 807 648 841 674
rect 807 640 841 648
rect 807 580 841 602
rect 807 568 841 580
rect 807 512 841 530
rect 807 496 841 512
rect 807 444 841 458
rect 807 424 841 444
rect 807 376 841 386
rect 807 352 841 376
rect 807 308 841 314
rect 807 280 841 308
rect 807 240 841 242
rect 807 208 841 240
rect 807 138 841 170
rect 807 136 841 138
rect 942 1464 976 1466
rect 942 1432 976 1464
rect 942 1362 976 1394
rect 942 1360 976 1362
rect 942 1294 976 1322
rect 942 1288 976 1294
rect 942 1226 976 1250
rect 942 1216 976 1226
rect 942 1158 976 1178
rect 942 1144 976 1158
rect 942 1090 976 1106
rect 942 1072 976 1090
rect 942 1022 976 1034
rect 942 1000 976 1022
rect 942 954 976 962
rect 942 928 976 954
rect 942 886 976 890
rect 942 856 976 886
rect 942 784 976 818
rect 942 716 976 746
rect 942 712 976 716
rect 942 648 976 674
rect 942 640 976 648
rect 942 580 976 602
rect 942 568 976 580
rect 942 512 976 530
rect 942 496 976 512
rect 942 444 976 458
rect 942 424 976 444
rect 942 376 976 386
rect 942 352 976 376
rect 942 308 976 314
rect 942 280 976 308
rect 942 240 976 242
rect 942 208 976 240
rect 942 138 976 170
rect 942 136 976 138
rect 243 20 257 54
rect 257 20 277 54
rect 315 20 325 54
rect 325 20 349 54
rect 387 20 393 54
rect 393 20 421 54
rect 459 20 461 54
rect 461 20 493 54
rect 531 20 563 54
rect 563 20 565 54
rect 603 20 631 54
rect 631 20 637 54
rect 675 20 699 54
rect 699 20 709 54
rect 747 20 767 54
rect 767 20 781 54
<< metal1 >>
rect 231 1582 793 1602
rect 231 1548 243 1582
rect 277 1548 315 1582
rect 349 1548 387 1582
rect 421 1548 459 1582
rect 493 1548 531 1582
rect 565 1548 603 1582
rect 637 1548 675 1582
rect 709 1548 747 1582
rect 781 1548 793 1582
rect 231 1536 793 1548
rect 36 1466 94 1497
rect 36 1432 48 1466
rect 82 1432 94 1466
rect 36 1394 94 1432
rect 36 1360 48 1394
rect 82 1360 94 1394
rect 36 1322 94 1360
rect 36 1288 48 1322
rect 82 1288 94 1322
rect 36 1250 94 1288
rect 36 1216 48 1250
rect 82 1216 94 1250
rect 36 1178 94 1216
rect 36 1144 48 1178
rect 82 1144 94 1178
rect 36 1106 94 1144
rect 36 1072 48 1106
rect 82 1072 94 1106
rect 36 1034 94 1072
rect 36 1000 48 1034
rect 82 1000 94 1034
rect 36 962 94 1000
rect 36 928 48 962
rect 82 928 94 962
rect 36 890 94 928
rect 36 856 48 890
rect 82 856 94 890
rect 36 818 94 856
rect 36 784 48 818
rect 82 784 94 818
rect 36 746 94 784
rect 36 712 48 746
rect 82 712 94 746
rect 36 674 94 712
rect 36 640 48 674
rect 82 640 94 674
rect 36 602 94 640
rect 36 568 48 602
rect 82 568 94 602
rect 36 530 94 568
rect 36 496 48 530
rect 82 496 94 530
rect 36 458 94 496
rect 36 424 48 458
rect 82 424 94 458
rect 36 386 94 424
rect 36 352 48 386
rect 82 352 94 386
rect 36 314 94 352
rect 36 280 48 314
rect 82 280 94 314
rect 36 242 94 280
rect 36 208 48 242
rect 82 208 94 242
rect 36 170 94 208
rect 36 136 48 170
rect 82 136 94 170
rect 36 105 94 136
rect 174 1491 226 1497
rect 174 1432 183 1439
rect 217 1432 226 1439
rect 174 1427 226 1432
rect 174 1363 183 1375
rect 217 1363 226 1375
rect 174 1299 183 1311
rect 217 1299 226 1311
rect 174 1235 183 1247
rect 217 1235 226 1247
rect 174 1178 226 1183
rect 174 1144 183 1178
rect 217 1144 226 1178
rect 174 1106 226 1144
rect 174 1072 183 1106
rect 217 1072 226 1106
rect 174 1034 226 1072
rect 174 1000 183 1034
rect 217 1000 226 1034
rect 174 962 226 1000
rect 174 928 183 962
rect 217 928 226 962
rect 174 890 226 928
rect 174 856 183 890
rect 217 856 226 890
rect 174 818 226 856
rect 174 784 183 818
rect 217 784 226 818
rect 174 746 226 784
rect 174 712 183 746
rect 217 712 226 746
rect 174 674 226 712
rect 174 640 183 674
rect 217 640 226 674
rect 174 602 226 640
rect 174 568 183 602
rect 217 568 226 602
rect 174 530 226 568
rect 174 496 183 530
rect 217 496 226 530
rect 174 458 226 496
rect 174 424 183 458
rect 217 424 226 458
rect 174 419 226 424
rect 174 355 183 367
rect 217 355 226 367
rect 174 291 183 303
rect 217 291 226 303
rect 174 227 183 239
rect 217 227 226 239
rect 174 170 226 175
rect 174 163 183 170
rect 217 163 226 170
rect 174 105 226 111
rect 330 1466 382 1497
rect 330 1432 339 1466
rect 373 1432 382 1466
rect 330 1394 382 1432
rect 330 1360 339 1394
rect 373 1360 382 1394
rect 330 1322 382 1360
rect 330 1288 339 1322
rect 373 1288 382 1322
rect 330 1250 382 1288
rect 330 1216 339 1250
rect 373 1216 382 1250
rect 330 1178 382 1216
rect 330 1144 339 1178
rect 373 1144 382 1178
rect 330 1115 382 1144
rect 330 1051 382 1063
rect 330 987 382 999
rect 330 928 339 935
rect 373 928 382 935
rect 330 923 382 928
rect 330 859 339 871
rect 373 859 382 871
rect 330 795 339 807
rect 373 795 382 807
rect 330 731 339 743
rect 373 731 382 743
rect 330 674 382 679
rect 330 667 339 674
rect 373 667 382 674
rect 330 603 382 615
rect 330 539 382 551
rect 330 458 382 487
rect 330 424 339 458
rect 373 424 382 458
rect 330 386 382 424
rect 330 352 339 386
rect 373 352 382 386
rect 330 314 382 352
rect 330 280 339 314
rect 373 280 382 314
rect 330 242 382 280
rect 330 208 339 242
rect 373 208 382 242
rect 330 170 382 208
rect 330 136 339 170
rect 373 136 382 170
rect 330 105 382 136
rect 486 1491 538 1497
rect 486 1432 495 1439
rect 529 1432 538 1439
rect 486 1427 538 1432
rect 486 1363 495 1375
rect 529 1363 538 1375
rect 486 1299 495 1311
rect 529 1299 538 1311
rect 486 1235 495 1247
rect 529 1235 538 1247
rect 486 1178 538 1183
rect 486 1144 495 1178
rect 529 1144 538 1178
rect 486 1106 538 1144
rect 486 1072 495 1106
rect 529 1072 538 1106
rect 486 1034 538 1072
rect 486 1000 495 1034
rect 529 1000 538 1034
rect 486 962 538 1000
rect 486 928 495 962
rect 529 928 538 962
rect 486 890 538 928
rect 486 856 495 890
rect 529 856 538 890
rect 486 818 538 856
rect 486 784 495 818
rect 529 784 538 818
rect 486 746 538 784
rect 486 712 495 746
rect 529 712 538 746
rect 486 674 538 712
rect 486 640 495 674
rect 529 640 538 674
rect 486 602 538 640
rect 486 568 495 602
rect 529 568 538 602
rect 486 530 538 568
rect 486 496 495 530
rect 529 496 538 530
rect 486 458 538 496
rect 486 424 495 458
rect 529 424 538 458
rect 486 419 538 424
rect 486 355 495 367
rect 529 355 538 367
rect 486 291 495 303
rect 529 291 538 303
rect 486 227 495 239
rect 529 227 538 239
rect 486 170 538 175
rect 486 163 495 170
rect 529 163 538 170
rect 486 105 538 111
rect 642 1466 694 1497
rect 642 1432 651 1466
rect 685 1432 694 1466
rect 642 1394 694 1432
rect 642 1360 651 1394
rect 685 1360 694 1394
rect 642 1322 694 1360
rect 642 1288 651 1322
rect 685 1288 694 1322
rect 642 1250 694 1288
rect 642 1216 651 1250
rect 685 1216 694 1250
rect 642 1178 694 1216
rect 642 1144 651 1178
rect 685 1144 694 1178
rect 642 1115 694 1144
rect 642 1051 694 1063
rect 642 987 694 999
rect 642 928 651 935
rect 685 928 694 935
rect 642 923 694 928
rect 642 859 651 871
rect 685 859 694 871
rect 642 795 651 807
rect 685 795 694 807
rect 642 731 651 743
rect 685 731 694 743
rect 642 674 694 679
rect 642 667 651 674
rect 685 667 694 674
rect 642 603 694 615
rect 642 539 694 551
rect 642 458 694 487
rect 642 424 651 458
rect 685 424 694 458
rect 642 386 694 424
rect 642 352 651 386
rect 685 352 694 386
rect 642 314 694 352
rect 642 280 651 314
rect 685 280 694 314
rect 642 242 694 280
rect 642 208 651 242
rect 685 208 694 242
rect 642 170 694 208
rect 642 136 651 170
rect 685 136 694 170
rect 642 105 694 136
rect 798 1491 850 1497
rect 798 1432 807 1439
rect 841 1432 850 1439
rect 798 1427 850 1432
rect 798 1363 807 1375
rect 841 1363 850 1375
rect 798 1299 807 1311
rect 841 1299 850 1311
rect 798 1235 807 1247
rect 841 1235 850 1247
rect 798 1178 850 1183
rect 798 1144 807 1178
rect 841 1144 850 1178
rect 798 1106 850 1144
rect 798 1072 807 1106
rect 841 1072 850 1106
rect 798 1034 850 1072
rect 798 1000 807 1034
rect 841 1000 850 1034
rect 798 962 850 1000
rect 798 928 807 962
rect 841 928 850 962
rect 798 890 850 928
rect 798 856 807 890
rect 841 856 850 890
rect 798 818 850 856
rect 798 784 807 818
rect 841 784 850 818
rect 798 746 850 784
rect 798 712 807 746
rect 841 712 850 746
rect 798 674 850 712
rect 798 640 807 674
rect 841 640 850 674
rect 798 602 850 640
rect 798 568 807 602
rect 841 568 850 602
rect 798 530 850 568
rect 798 496 807 530
rect 841 496 850 530
rect 798 458 850 496
rect 798 424 807 458
rect 841 424 850 458
rect 798 419 850 424
rect 798 355 807 367
rect 841 355 850 367
rect 798 291 807 303
rect 841 291 850 303
rect 798 227 807 239
rect 841 227 850 239
rect 798 170 850 175
rect 798 163 807 170
rect 841 163 850 170
rect 798 105 850 111
rect 930 1466 988 1497
rect 930 1432 942 1466
rect 976 1432 988 1466
rect 930 1394 988 1432
rect 930 1360 942 1394
rect 976 1360 988 1394
rect 930 1322 988 1360
rect 930 1288 942 1322
rect 976 1288 988 1322
rect 930 1250 988 1288
rect 930 1216 942 1250
rect 976 1216 988 1250
rect 930 1178 988 1216
rect 930 1144 942 1178
rect 976 1144 988 1178
rect 930 1106 988 1144
rect 930 1072 942 1106
rect 976 1072 988 1106
rect 930 1034 988 1072
rect 930 1000 942 1034
rect 976 1000 988 1034
rect 930 962 988 1000
rect 930 928 942 962
rect 976 928 988 962
rect 930 890 988 928
rect 930 856 942 890
rect 976 856 988 890
rect 930 818 988 856
rect 930 784 942 818
rect 976 784 988 818
rect 930 746 988 784
rect 930 712 942 746
rect 976 712 988 746
rect 930 674 988 712
rect 930 640 942 674
rect 976 640 988 674
rect 930 602 988 640
rect 930 568 942 602
rect 976 568 988 602
rect 930 530 988 568
rect 930 496 942 530
rect 976 496 988 530
rect 930 458 988 496
rect 930 424 942 458
rect 976 424 988 458
rect 930 386 988 424
rect 930 352 942 386
rect 976 352 988 386
rect 930 314 988 352
rect 930 280 942 314
rect 976 280 988 314
rect 930 242 988 280
rect 930 208 942 242
rect 976 208 988 242
rect 930 170 988 208
rect 930 136 942 170
rect 976 136 988 170
rect 930 105 988 136
rect 231 54 793 66
rect 231 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 531 54
rect 565 20 603 54
rect 637 20 675 54
rect 709 20 747 54
rect 781 20 793 54
rect 231 0 793 20
<< via1 >>
rect 174 1466 226 1491
rect 174 1439 183 1466
rect 183 1439 217 1466
rect 217 1439 226 1466
rect 174 1394 226 1427
rect 174 1375 183 1394
rect 183 1375 217 1394
rect 217 1375 226 1394
rect 174 1360 183 1363
rect 183 1360 217 1363
rect 217 1360 226 1363
rect 174 1322 226 1360
rect 174 1311 183 1322
rect 183 1311 217 1322
rect 217 1311 226 1322
rect 174 1288 183 1299
rect 183 1288 217 1299
rect 217 1288 226 1299
rect 174 1250 226 1288
rect 174 1247 183 1250
rect 183 1247 217 1250
rect 217 1247 226 1250
rect 174 1216 183 1235
rect 183 1216 217 1235
rect 217 1216 226 1235
rect 174 1183 226 1216
rect 174 386 226 419
rect 174 367 183 386
rect 183 367 217 386
rect 217 367 226 386
rect 174 352 183 355
rect 183 352 217 355
rect 217 352 226 355
rect 174 314 226 352
rect 174 303 183 314
rect 183 303 217 314
rect 217 303 226 314
rect 174 280 183 291
rect 183 280 217 291
rect 217 280 226 291
rect 174 242 226 280
rect 174 239 183 242
rect 183 239 217 242
rect 217 239 226 242
rect 174 208 183 227
rect 183 208 217 227
rect 217 208 226 227
rect 174 175 226 208
rect 174 136 183 163
rect 183 136 217 163
rect 217 136 226 163
rect 174 111 226 136
rect 330 1106 382 1115
rect 330 1072 339 1106
rect 339 1072 373 1106
rect 373 1072 382 1106
rect 330 1063 382 1072
rect 330 1034 382 1051
rect 330 1000 339 1034
rect 339 1000 373 1034
rect 373 1000 382 1034
rect 330 999 382 1000
rect 330 962 382 987
rect 330 935 339 962
rect 339 935 373 962
rect 373 935 382 962
rect 330 890 382 923
rect 330 871 339 890
rect 339 871 373 890
rect 373 871 382 890
rect 330 856 339 859
rect 339 856 373 859
rect 373 856 382 859
rect 330 818 382 856
rect 330 807 339 818
rect 339 807 373 818
rect 373 807 382 818
rect 330 784 339 795
rect 339 784 373 795
rect 373 784 382 795
rect 330 746 382 784
rect 330 743 339 746
rect 339 743 373 746
rect 373 743 382 746
rect 330 712 339 731
rect 339 712 373 731
rect 373 712 382 731
rect 330 679 382 712
rect 330 640 339 667
rect 339 640 373 667
rect 373 640 382 667
rect 330 615 382 640
rect 330 602 382 603
rect 330 568 339 602
rect 339 568 373 602
rect 373 568 382 602
rect 330 551 382 568
rect 330 530 382 539
rect 330 496 339 530
rect 339 496 373 530
rect 373 496 382 530
rect 330 487 382 496
rect 486 1466 538 1491
rect 486 1439 495 1466
rect 495 1439 529 1466
rect 529 1439 538 1466
rect 486 1394 538 1427
rect 486 1375 495 1394
rect 495 1375 529 1394
rect 529 1375 538 1394
rect 486 1360 495 1363
rect 495 1360 529 1363
rect 529 1360 538 1363
rect 486 1322 538 1360
rect 486 1311 495 1322
rect 495 1311 529 1322
rect 529 1311 538 1322
rect 486 1288 495 1299
rect 495 1288 529 1299
rect 529 1288 538 1299
rect 486 1250 538 1288
rect 486 1247 495 1250
rect 495 1247 529 1250
rect 529 1247 538 1250
rect 486 1216 495 1235
rect 495 1216 529 1235
rect 529 1216 538 1235
rect 486 1183 538 1216
rect 486 386 538 419
rect 486 367 495 386
rect 495 367 529 386
rect 529 367 538 386
rect 486 352 495 355
rect 495 352 529 355
rect 529 352 538 355
rect 486 314 538 352
rect 486 303 495 314
rect 495 303 529 314
rect 529 303 538 314
rect 486 280 495 291
rect 495 280 529 291
rect 529 280 538 291
rect 486 242 538 280
rect 486 239 495 242
rect 495 239 529 242
rect 529 239 538 242
rect 486 208 495 227
rect 495 208 529 227
rect 529 208 538 227
rect 486 175 538 208
rect 486 136 495 163
rect 495 136 529 163
rect 529 136 538 163
rect 486 111 538 136
rect 642 1106 694 1115
rect 642 1072 651 1106
rect 651 1072 685 1106
rect 685 1072 694 1106
rect 642 1063 694 1072
rect 642 1034 694 1051
rect 642 1000 651 1034
rect 651 1000 685 1034
rect 685 1000 694 1034
rect 642 999 694 1000
rect 642 962 694 987
rect 642 935 651 962
rect 651 935 685 962
rect 685 935 694 962
rect 642 890 694 923
rect 642 871 651 890
rect 651 871 685 890
rect 685 871 694 890
rect 642 856 651 859
rect 651 856 685 859
rect 685 856 694 859
rect 642 818 694 856
rect 642 807 651 818
rect 651 807 685 818
rect 685 807 694 818
rect 642 784 651 795
rect 651 784 685 795
rect 685 784 694 795
rect 642 746 694 784
rect 642 743 651 746
rect 651 743 685 746
rect 685 743 694 746
rect 642 712 651 731
rect 651 712 685 731
rect 685 712 694 731
rect 642 679 694 712
rect 642 640 651 667
rect 651 640 685 667
rect 685 640 694 667
rect 642 615 694 640
rect 642 602 694 603
rect 642 568 651 602
rect 651 568 685 602
rect 685 568 694 602
rect 642 551 694 568
rect 642 530 694 539
rect 642 496 651 530
rect 651 496 685 530
rect 685 496 694 530
rect 642 487 694 496
rect 798 1466 850 1491
rect 798 1439 807 1466
rect 807 1439 841 1466
rect 841 1439 850 1466
rect 798 1394 850 1427
rect 798 1375 807 1394
rect 807 1375 841 1394
rect 841 1375 850 1394
rect 798 1360 807 1363
rect 807 1360 841 1363
rect 841 1360 850 1363
rect 798 1322 850 1360
rect 798 1311 807 1322
rect 807 1311 841 1322
rect 841 1311 850 1322
rect 798 1288 807 1299
rect 807 1288 841 1299
rect 841 1288 850 1299
rect 798 1250 850 1288
rect 798 1247 807 1250
rect 807 1247 841 1250
rect 841 1247 850 1250
rect 798 1216 807 1235
rect 807 1216 841 1235
rect 841 1216 850 1235
rect 798 1183 850 1216
rect 798 386 850 419
rect 798 367 807 386
rect 807 367 841 386
rect 841 367 850 386
rect 798 352 807 355
rect 807 352 841 355
rect 841 352 850 355
rect 798 314 850 352
rect 798 303 807 314
rect 807 303 841 314
rect 841 303 850 314
rect 798 280 807 291
rect 807 280 841 291
rect 841 280 850 291
rect 798 242 850 280
rect 798 239 807 242
rect 807 239 841 242
rect 841 239 850 242
rect 798 208 807 227
rect 807 208 841 227
rect 841 208 850 227
rect 798 175 850 208
rect 798 136 807 163
rect 807 136 841 163
rect 841 136 850 163
rect 798 111 850 136
<< metal2 >>
rect 10 1491 1014 1497
rect 10 1439 174 1491
rect 226 1439 486 1491
rect 538 1439 798 1491
rect 850 1439 1014 1491
rect 10 1427 1014 1439
rect 10 1375 174 1427
rect 226 1375 486 1427
rect 538 1375 798 1427
rect 850 1375 1014 1427
rect 10 1363 1014 1375
rect 10 1311 174 1363
rect 226 1311 486 1363
rect 538 1311 798 1363
rect 850 1311 1014 1363
rect 10 1299 1014 1311
rect 10 1247 174 1299
rect 226 1247 486 1299
rect 538 1247 798 1299
rect 850 1247 1014 1299
rect 10 1235 1014 1247
rect 10 1183 174 1235
rect 226 1183 486 1235
rect 538 1183 798 1235
rect 850 1183 1014 1235
rect 10 1177 1014 1183
rect 10 1115 1014 1121
rect 10 1063 330 1115
rect 382 1063 642 1115
rect 694 1063 1014 1115
rect 10 1051 1014 1063
rect 10 999 330 1051
rect 382 999 642 1051
rect 694 999 1014 1051
rect 10 987 1014 999
rect 10 935 330 987
rect 382 935 642 987
rect 694 935 1014 987
rect 10 923 1014 935
rect 10 871 330 923
rect 382 871 642 923
rect 694 871 1014 923
rect 10 859 1014 871
rect 10 807 330 859
rect 382 807 642 859
rect 694 807 1014 859
rect 10 795 1014 807
rect 10 743 330 795
rect 382 743 642 795
rect 694 743 1014 795
rect 10 731 1014 743
rect 10 679 330 731
rect 382 679 642 731
rect 694 679 1014 731
rect 10 667 1014 679
rect 10 615 330 667
rect 382 615 642 667
rect 694 615 1014 667
rect 10 603 1014 615
rect 10 551 330 603
rect 382 551 642 603
rect 694 551 1014 603
rect 10 539 1014 551
rect 10 487 330 539
rect 382 487 642 539
rect 694 487 1014 539
rect 10 481 1014 487
rect 10 419 1014 425
rect 10 367 174 419
rect 226 367 486 419
rect 538 367 798 419
rect 850 367 1014 419
rect 10 355 1014 367
rect 10 303 174 355
rect 226 303 486 355
rect 538 303 798 355
rect 850 303 1014 355
rect 10 291 1014 303
rect 10 239 174 291
rect 226 239 486 291
rect 538 239 798 291
rect 850 239 1014 291
rect 10 227 1014 239
rect 10 175 174 227
rect 226 175 486 227
rect 538 175 798 227
rect 850 175 1014 227
rect 10 163 1014 175
rect 10 111 174 163
rect 226 111 486 163
rect 538 111 798 163
rect 850 111 1014 163
rect 10 105 1014 111
<< labels >>
flabel comment s 824 801 824 801 0 FreeSans 300 0 0 0 S
flabel comment s 668 801 668 801 0 FreeSans 300 0 0 0 S
flabel comment s 668 801 668 801 0 FreeSans 300 0 0 0 D
flabel comment s 512 801 512 801 0 FreeSans 300 0 0 0 S
flabel comment s 512 801 512 801 0 FreeSans 300 0 0 0 S
flabel comment s 356 801 356 801 0 FreeSans 300 0 0 0 S
flabel comment s 356 801 356 801 0 FreeSans 300 0 0 0 D
flabel comment s 200 801 200 801 0 FreeSans 300 0 0 0 S
flabel comment s 200 801 200 801 0 FreeSans 300 0 0 0 S
flabel metal1 s 449 1551 569 1584 0 FreeSans 200 0 0 0 GATE
flabel metal1 s 441 15 575 54 0 FreeSans 200 0 0 0 GATE
flabel metal1 s 53 1007 83 1264 0 FreeSans 200 90 0 0 SUBSTRATE
flabel metal1 s 944 1028 968 1270 0 FreeSans 200 90 0 0 SUBSTRATE
flabel metal2 s 107 683 148 919 0 FreeSans 200 90 0 0 DRAIN
flabel metal2 s 50 1259 86 1420 0 FreeSans 200 90 0 0 SOURCE
flabel metal2 s 47 153 89 349 0 FreeSans 200 90 0 0 SOURCE
<< properties >>
string GDS_END 4348170
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4318450
<< end >>
