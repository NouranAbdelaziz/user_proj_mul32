magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect 0 0 604 806
<< pmoslvt >>
rect 204 102 274 704
rect 330 102 400 704
<< pdiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 274 692 330 704
rect 274 658 285 692
rect 319 658 330 692
rect 274 624 330 658
rect 274 590 285 624
rect 319 590 330 624
rect 274 556 330 590
rect 274 522 285 556
rect 319 522 330 556
rect 274 488 330 522
rect 274 454 285 488
rect 319 454 330 488
rect 274 420 330 454
rect 274 386 285 420
rect 319 386 330 420
rect 274 352 330 386
rect 274 318 285 352
rect 319 318 330 352
rect 274 284 330 318
rect 274 250 285 284
rect 319 250 330 284
rect 274 216 330 250
rect 274 182 285 216
rect 319 182 330 216
rect 274 148 330 182
rect 274 114 285 148
rect 319 114 330 148
rect 274 102 330 114
rect 400 692 456 704
rect 400 658 411 692
rect 445 658 456 692
rect 400 624 456 658
rect 400 590 411 624
rect 445 590 456 624
rect 400 556 456 590
rect 400 522 411 556
rect 445 522 456 556
rect 400 488 456 522
rect 400 454 411 488
rect 445 454 456 488
rect 400 420 456 454
rect 400 386 411 420
rect 445 386 456 420
rect 400 352 456 386
rect 400 318 411 352
rect 445 318 456 352
rect 400 284 456 318
rect 400 250 411 284
rect 445 250 456 284
rect 400 216 456 250
rect 400 182 411 216
rect 445 182 456 216
rect 400 148 456 182
rect 400 114 411 148
rect 445 114 456 148
rect 400 102 456 114
<< pdiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 285 658 319 692
rect 285 590 319 624
rect 285 522 319 556
rect 285 454 319 488
rect 285 386 319 420
rect 285 318 319 352
rect 285 250 319 284
rect 285 182 319 216
rect 285 114 319 148
rect 411 658 445 692
rect 411 590 445 624
rect 411 522 445 556
rect 411 454 445 488
rect 411 386 445 420
rect 411 318 445 352
rect 411 250 445 284
rect 411 182 445 216
rect 411 114 445 148
<< nsubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 510 658 568 704
rect 510 624 522 658
rect 556 624 568 658
rect 510 590 568 624
rect 510 556 522 590
rect 556 556 568 590
rect 510 522 568 556
rect 510 488 522 522
rect 556 488 568 522
rect 510 454 568 488
rect 510 420 522 454
rect 556 420 568 454
rect 510 386 568 420
rect 510 352 522 386
rect 556 352 568 386
rect 510 318 568 352
rect 510 284 522 318
rect 556 284 568 318
rect 510 250 568 284
rect 510 216 522 250
rect 556 216 568 250
rect 510 182 568 216
rect 510 148 522 182
rect 556 148 568 182
rect 510 102 568 148
<< nsubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 522 624 556 658
rect 522 556 556 590
rect 522 488 556 522
rect 522 420 556 454
rect 522 352 556 386
rect 522 284 556 318
rect 522 216 556 250
rect 522 148 556 182
<< poly >>
rect 165 786 439 806
rect 165 752 183 786
rect 217 752 251 786
rect 285 752 319 786
rect 353 752 387 786
rect 421 752 439 786
rect 165 736 439 752
rect 204 704 274 736
rect 330 704 400 736
rect 204 70 274 102
rect 330 70 400 102
rect 165 54 439 70
rect 165 20 183 54
rect 217 20 251 54
rect 285 20 319 54
rect 353 20 387 54
rect 421 20 439 54
rect 165 0 439 20
<< polycont >>
rect 183 752 217 786
rect 251 752 285 786
rect 319 752 353 786
rect 387 752 421 786
rect 183 20 217 54
rect 251 20 285 54
rect 319 20 353 54
rect 387 20 421 54
<< locali >>
rect 165 752 177 786
rect 217 752 249 786
rect 285 752 319 786
rect 355 752 387 786
rect 427 752 439 786
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 285 692 319 708
rect 285 624 319 638
rect 285 556 319 566
rect 285 488 319 494
rect 285 420 319 422
rect 285 384 319 386
rect 285 312 319 318
rect 285 240 319 250
rect 285 168 319 182
rect 285 98 319 114
rect 411 692 445 708
rect 411 624 445 638
rect 411 556 445 566
rect 411 488 445 494
rect 411 420 445 422
rect 411 384 445 386
rect 411 312 445 318
rect 411 240 445 250
rect 411 168 445 182
rect 522 672 556 674
rect 522 600 556 624
rect 522 528 556 556
rect 522 456 556 488
rect 522 386 556 420
rect 522 318 556 350
rect 522 250 556 278
rect 522 182 556 206
rect 522 132 556 134
rect 411 98 445 114
rect 165 20 177 54
rect 217 20 249 54
rect 285 20 319 54
rect 355 20 387 54
rect 427 20 439 54
<< viali >>
rect 177 752 183 786
rect 183 752 211 786
rect 249 752 251 786
rect 251 752 283 786
rect 321 752 353 786
rect 353 752 355 786
rect 393 752 421 786
rect 421 752 427 786
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 285 658 319 672
rect 285 638 319 658
rect 285 590 319 600
rect 285 566 319 590
rect 285 522 319 528
rect 285 494 319 522
rect 285 454 319 456
rect 285 422 319 454
rect 285 352 319 384
rect 285 350 319 352
rect 285 284 319 312
rect 285 278 319 284
rect 285 216 319 240
rect 285 206 319 216
rect 285 148 319 168
rect 285 134 319 148
rect 411 658 445 672
rect 411 638 445 658
rect 411 590 445 600
rect 411 566 445 590
rect 411 522 445 528
rect 411 494 445 522
rect 411 454 445 456
rect 411 422 445 454
rect 411 352 445 384
rect 411 350 445 352
rect 411 284 445 312
rect 411 278 445 284
rect 411 216 445 240
rect 411 206 445 216
rect 411 148 445 168
rect 411 134 445 148
rect 522 658 556 672
rect 522 638 556 658
rect 522 590 556 600
rect 522 566 556 590
rect 522 522 556 528
rect 522 494 556 522
rect 522 454 556 456
rect 522 422 556 454
rect 522 352 556 384
rect 522 350 556 352
rect 522 284 556 312
rect 522 278 556 284
rect 522 216 556 240
rect 522 206 556 216
rect 522 148 556 168
rect 522 134 556 148
rect 177 20 183 54
rect 183 20 211 54
rect 249 20 251 54
rect 251 20 283 54
rect 321 20 353 54
rect 353 20 355 54
rect 393 20 421 54
rect 421 20 427 54
<< metal1 >>
rect 165 786 439 806
rect 165 752 177 786
rect 211 752 249 786
rect 283 752 321 786
rect 355 752 393 786
rect 427 752 439 786
rect 165 740 439 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 276 678 328 684
rect 276 614 328 626
rect 276 550 328 562
rect 276 494 285 498
rect 319 494 328 498
rect 276 486 328 494
rect 276 422 285 434
rect 319 422 328 434
rect 276 384 328 422
rect 276 350 285 384
rect 319 350 328 384
rect 276 312 328 350
rect 276 278 285 312
rect 319 278 328 312
rect 276 240 328 278
rect 276 206 285 240
rect 319 206 328 240
rect 276 168 328 206
rect 276 134 285 168
rect 319 134 328 168
rect 276 122 328 134
rect 402 672 454 684
rect 402 638 411 672
rect 445 638 454 672
rect 402 600 454 638
rect 402 566 411 600
rect 445 566 454 600
rect 402 528 454 566
rect 402 494 411 528
rect 445 494 454 528
rect 402 456 454 494
rect 402 422 411 456
rect 445 422 454 456
rect 402 384 454 422
rect 402 372 411 384
rect 445 372 454 384
rect 402 312 454 320
rect 402 308 411 312
rect 445 308 454 312
rect 402 244 454 256
rect 402 180 454 192
rect 402 122 454 128
rect 510 672 568 684
rect 510 638 522 672
rect 556 638 568 672
rect 510 600 568 638
rect 510 566 522 600
rect 556 566 568 600
rect 510 528 568 566
rect 510 494 522 528
rect 556 494 568 528
rect 510 456 568 494
rect 510 422 522 456
rect 556 422 568 456
rect 510 384 568 422
rect 510 350 522 384
rect 556 350 568 384
rect 510 312 568 350
rect 510 278 522 312
rect 556 278 568 312
rect 510 240 568 278
rect 510 206 522 240
rect 556 206 568 240
rect 510 168 568 206
rect 510 134 522 168
rect 556 134 568 168
rect 510 122 568 134
rect 165 54 439 66
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 439 54
rect 165 0 439 20
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 276 672 328 678
rect 276 638 285 672
rect 285 638 319 672
rect 319 638 328 672
rect 276 626 328 638
rect 276 600 328 614
rect 276 566 285 600
rect 285 566 319 600
rect 319 566 328 600
rect 276 562 328 566
rect 276 528 328 550
rect 276 498 285 528
rect 285 498 319 528
rect 319 498 328 528
rect 276 456 328 486
rect 276 434 285 456
rect 285 434 319 456
rect 319 434 328 456
rect 402 350 411 372
rect 411 350 445 372
rect 445 350 454 372
rect 402 320 454 350
rect 402 278 411 308
rect 411 278 445 308
rect 445 278 454 308
rect 402 256 454 278
rect 402 240 454 244
rect 402 206 411 240
rect 411 206 445 240
rect 445 206 454 240
rect 402 192 454 206
rect 402 168 454 180
rect 402 134 411 168
rect 411 134 445 168
rect 445 134 454 168
rect 402 128 454 134
<< metal2 >>
rect 10 678 594 684
rect 10 626 276 678
rect 328 626 594 678
rect 10 614 594 626
rect 10 562 276 614
rect 328 562 594 614
rect 10 550 594 562
rect 10 498 276 550
rect 328 498 594 550
rect 10 486 594 498
rect 10 434 276 486
rect 328 434 594 486
rect 10 428 594 434
rect 10 372 594 378
rect 10 320 150 372
rect 202 320 402 372
rect 454 320 594 372
rect 10 308 594 320
rect 10 256 150 308
rect 202 256 402 308
rect 454 256 594 308
rect 10 244 594 256
rect 10 192 150 244
rect 202 192 402 244
rect 454 192 594 244
rect 10 180 594 192
rect 10 128 150 180
rect 202 128 402 180
rect 454 128 594 180
rect 10 122 594 128
<< labels >>
flabel metal2 s 10 122 30 378 7 FreeSans 300 180 0 0 SOURCE
flabel metal2 s 10 428 30 684 7 FreeSans 300 180 0 0 DRAIN
flabel metal1 s 165 0 439 66 0 FreeSans 300 0 0 0 GATE
flabel metal1 s 165 740 439 806 0 FreeSans 300 0 0 0 GATE
flabel metal1 s 510 122 568 138 3 FreeSans 300 90 0 0 BULK
flabel metal1 s 36 122 94 138 3 FreeSans 300 90 0 0 BULK
<< properties >>
string GDS_END 9849686
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9838578
<< end >>
