/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.ref/sky130_sram_macros/spice/sky130_sram_1kbyte_1rw1r_8x1024_8.spice