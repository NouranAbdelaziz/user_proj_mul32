/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/capacitors/sky130_fd_pr__model__cap_var.model.spice