* NGSPICE file created from sky130_ef_sc_hd__fill_4.ext - technology: sky130B

.subckt sky130_ef_sc_hd__fill_4
.ends

