/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/correl2.spice