/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8_mvt.pm3.spice