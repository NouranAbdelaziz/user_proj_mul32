/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/parameters/slow.spice