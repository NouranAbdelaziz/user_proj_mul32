magic
tech sky130A
magscale 1 2
timestamp 1685891715
<< nwell >>
rect 1066 349509 558846 349830
rect 1066 348421 558846 348987
rect 1066 347333 558846 347899
rect 1066 346245 558846 346811
rect 1066 345157 558846 345723
rect 1066 344069 558846 344635
rect 1066 342981 558846 343547
rect 1066 341893 558846 342459
rect 1066 340805 558846 341371
rect 1066 339717 558846 340283
rect 1066 338629 558846 339195
rect 1066 337541 558846 338107
rect 1066 336453 558846 337019
rect 1066 335365 558846 335931
rect 1066 334277 558846 334843
rect 1066 333189 558846 333755
rect 1066 332101 558846 332667
rect 1066 331013 558846 331579
rect 1066 329925 558846 330491
rect 1066 328837 558846 329403
rect 1066 327749 558846 328315
rect 1066 326661 558846 327227
rect 1066 325573 558846 326139
rect 1066 324485 558846 325051
rect 1066 323397 558846 323963
rect 1066 322309 558846 322875
rect 1066 321221 558846 321787
rect 1066 320133 558846 320699
rect 1066 319045 558846 319611
rect 1066 317957 558846 318523
rect 1066 316869 558846 317435
rect 1066 315781 558846 316347
rect 1066 314693 558846 315259
rect 1066 313605 558846 314171
rect 1066 312517 558846 313083
rect 1066 311429 558846 311995
rect 1066 310341 558846 310907
rect 1066 309253 558846 309819
rect 1066 308165 558846 308731
rect 1066 307077 558846 307643
rect 1066 305989 558846 306555
rect 1066 304901 558846 305467
rect 1066 303813 558846 304379
rect 1066 302725 558846 303291
rect 1066 301637 558846 302203
rect 1066 300549 558846 301115
rect 1066 299461 558846 300027
rect 1066 298373 558846 298939
rect 1066 297285 558846 297851
rect 1066 296197 558846 296763
rect 1066 295109 558846 295675
rect 1066 294021 558846 294587
rect 1066 292933 558846 293499
rect 1066 291845 558846 292411
rect 1066 290757 558846 291323
rect 1066 289669 558846 290235
rect 1066 288581 558846 289147
rect 1066 287493 558846 288059
rect 1066 286405 558846 286971
rect 1066 285317 558846 285883
rect 1066 284229 558846 284795
rect 1066 283141 558846 283707
rect 1066 282053 558846 282619
rect 1066 280965 558846 281531
rect 1066 279877 558846 280443
rect 1066 278789 558846 279355
rect 1066 277701 558846 278267
rect 1066 276613 558846 277179
rect 1066 275525 558846 276091
rect 1066 274437 558846 275003
rect 1066 273349 558846 273915
rect 1066 272261 558846 272827
rect 1066 271173 558846 271739
rect 1066 270085 558846 270651
rect 1066 268997 558846 269563
rect 1066 267909 558846 268475
rect 1066 266821 558846 267387
rect 1066 265733 558846 266299
rect 1066 264645 558846 265211
rect 1066 263557 558846 264123
rect 1066 262469 558846 263035
rect 1066 261381 558846 261947
rect 1066 260293 558846 260859
rect 1066 259205 558846 259771
rect 1066 258117 558846 258683
rect 1066 257029 558846 257595
rect 1066 255941 558846 256507
rect 1066 254853 558846 255419
rect 1066 253765 558846 254331
rect 1066 252677 558846 253243
rect 1066 251589 558846 252155
rect 1066 250501 558846 251067
rect 1066 249413 558846 249979
rect 1066 248325 558846 248891
rect 1066 247237 558846 247803
rect 1066 246149 558846 246715
rect 1066 245061 558846 245627
rect 1066 243973 558846 244539
rect 1066 242885 558846 243451
rect 1066 241797 558846 242363
rect 1066 240709 558846 241275
rect 1066 239621 558846 240187
rect 1066 238533 558846 239099
rect 1066 237445 558846 238011
rect 1066 236357 558846 236923
rect 1066 235269 558846 235835
rect 1066 234181 558846 234747
rect 1066 233093 558846 233659
rect 1066 232005 558846 232571
rect 1066 230917 558846 231483
rect 1066 229829 558846 230395
rect 1066 228741 558846 229307
rect 1066 227653 558846 228219
rect 1066 226565 558846 227131
rect 1066 225477 558846 226043
rect 1066 224389 558846 224955
rect 1066 223301 558846 223867
rect 1066 222213 558846 222779
rect 1066 221125 558846 221691
rect 1066 220037 558846 220603
rect 1066 218949 558846 219515
rect 1066 217861 558846 218427
rect 1066 216773 558846 217339
rect 1066 215685 558846 216251
rect 1066 214597 558846 215163
rect 1066 213509 558846 214075
rect 1066 212421 558846 212987
rect 1066 211333 558846 211899
rect 1066 210245 558846 210811
rect 1066 209157 558846 209723
rect 1066 208069 558846 208635
rect 1066 206981 558846 207547
rect 1066 205893 558846 206459
rect 1066 204805 558846 205371
rect 1066 203717 558846 204283
rect 1066 202629 558846 203195
rect 1066 201541 558846 202107
rect 1066 200453 558846 201019
rect 1066 199365 558846 199931
rect 1066 198277 558846 198843
rect 1066 197189 558846 197755
rect 1066 196101 558846 196667
rect 1066 195013 558846 195579
rect 1066 193925 558846 194491
rect 1066 192837 558846 193403
rect 1066 191749 558846 192315
rect 1066 190661 558846 191227
rect 1066 189573 558846 190139
rect 1066 188485 558846 189051
rect 1066 187397 558846 187963
rect 1066 186309 558846 186875
rect 1066 185221 558846 185787
rect 1066 184133 558846 184699
rect 1066 183045 558846 183611
rect 1066 181957 558846 182523
rect 1066 180869 558846 181435
rect 1066 179781 558846 180347
rect 1066 178693 558846 179259
rect 1066 177605 558846 178171
rect 1066 176517 558846 177083
rect 1066 175429 558846 175995
rect 1066 174341 558846 174907
rect 1066 173253 558846 173819
rect 1066 172165 558846 172731
rect 1066 171077 558846 171643
rect 1066 169989 558846 170555
rect 1066 168901 558846 169467
rect 1066 167813 558846 168379
rect 1066 166725 558846 167291
rect 1066 165637 558846 166203
rect 1066 164549 558846 165115
rect 1066 163461 558846 164027
rect 1066 162373 558846 162939
rect 1066 161285 558846 161851
rect 1066 160197 558846 160763
rect 1066 159109 558846 159675
rect 1066 158021 558846 158587
rect 1066 156933 558846 157499
rect 1066 155845 558846 156411
rect 1066 154757 558846 155323
rect 1066 153669 558846 154235
rect 1066 152581 558846 153147
rect 1066 151493 558846 152059
rect 1066 150405 558846 150971
rect 1066 149317 558846 149883
rect 1066 148229 558846 148795
rect 1066 147141 558846 147707
rect 1066 146053 558846 146619
rect 1066 144965 558846 145531
rect 1066 143877 558846 144443
rect 1066 142789 558846 143355
rect 1066 141701 558846 142267
rect 1066 140613 558846 141179
rect 1066 139525 558846 140091
rect 1066 138437 558846 139003
rect 1066 137349 558846 137915
rect 1066 136261 558846 136827
rect 1066 135173 558846 135739
rect 1066 134085 558846 134651
rect 1066 132997 558846 133563
rect 1066 131909 558846 132475
rect 1066 130821 558846 131387
rect 1066 129733 558846 130299
rect 1066 128645 558846 129211
rect 1066 127557 558846 128123
rect 1066 126469 558846 127035
rect 1066 125381 558846 125947
rect 1066 124293 558846 124859
rect 1066 123205 558846 123771
rect 1066 122117 558846 122683
rect 1066 121029 558846 121595
rect 1066 119941 558846 120507
rect 1066 118853 558846 119419
rect 1066 117765 558846 118331
rect 1066 116677 558846 117243
rect 1066 115589 558846 116155
rect 1066 114501 558846 115067
rect 1066 113413 558846 113979
rect 1066 112325 558846 112891
rect 1066 111237 558846 111803
rect 1066 110149 558846 110715
rect 1066 109061 558846 109627
rect 1066 107973 558846 108539
rect 1066 106885 558846 107451
rect 1066 105797 558846 106363
rect 1066 104709 558846 105275
rect 1066 103621 558846 104187
rect 1066 102533 558846 103099
rect 1066 101445 558846 102011
rect 1066 100357 558846 100923
rect 1066 99269 558846 99835
rect 1066 98181 558846 98747
rect 1066 97093 558846 97659
rect 1066 96005 558846 96571
rect 1066 94917 558846 95483
rect 1066 93829 558846 94395
rect 1066 92741 558846 93307
rect 1066 91653 558846 92219
rect 1066 90565 558846 91131
rect 1066 89477 558846 90043
rect 1066 88389 558846 88955
rect 1066 87301 558846 87867
rect 1066 86213 558846 86779
rect 1066 85125 558846 85691
rect 1066 84037 558846 84603
rect 1066 82949 558846 83515
rect 1066 81861 558846 82427
rect 1066 80773 558846 81339
rect 1066 79685 558846 80251
rect 1066 78597 558846 79163
rect 1066 77509 558846 78075
rect 1066 76421 558846 76987
rect 1066 75333 558846 75899
rect 1066 74245 558846 74811
rect 1066 73157 558846 73723
rect 1066 72069 558846 72635
rect 1066 70981 558846 71547
rect 1066 69893 558846 70459
rect 1066 68805 558846 69371
rect 1066 67717 558846 68283
rect 1066 66629 558846 67195
rect 1066 65541 558846 66107
rect 1066 64453 558846 65019
rect 1066 63365 558846 63931
rect 1066 62277 558846 62843
rect 1066 61189 558846 61755
rect 1066 60101 558846 60667
rect 1066 59013 558846 59579
rect 1066 57925 558846 58491
rect 1066 56837 558846 57403
rect 1066 55749 558846 56315
rect 1066 54661 558846 55227
rect 1066 53573 558846 54139
rect 1066 52485 558846 53051
rect 1066 51397 558846 51963
rect 1066 50309 558846 50875
rect 1066 49221 558846 49787
rect 1066 48133 558846 48699
rect 1066 47045 558846 47611
rect 1066 45957 558846 46523
rect 1066 44869 558846 45435
rect 1066 43781 558846 44347
rect 1066 42693 558846 43259
rect 1066 41605 558846 42171
rect 1066 40517 558846 41083
rect 1066 39429 558846 39995
rect 1066 38341 558846 38907
rect 1066 37253 558846 37819
rect 1066 36165 558846 36731
rect 1066 35077 558846 35643
rect 1066 33989 558846 34555
rect 1066 32901 558846 33467
rect 1066 31813 558846 32379
rect 1066 30725 558846 31291
rect 1066 29637 558846 30203
rect 1066 28549 558846 29115
rect 1066 27461 558846 28027
rect 1066 26373 558846 26939
rect 1066 25285 558846 25851
rect 1066 24197 558846 24763
rect 1066 23109 558846 23675
rect 1066 22021 558846 22587
rect 1066 20933 558846 21499
rect 1066 19845 558846 20411
rect 1066 18757 558846 19323
rect 1066 17669 558846 18235
rect 1066 16581 558846 17147
rect 1066 15493 558846 16059
rect 1066 14405 558846 14971
rect 1066 13317 558846 13883
rect 1066 12229 558846 12795
rect 1066 11141 558846 11707
rect 1066 10053 558846 10619
rect 1066 8965 558846 9531
rect 1066 7877 558846 8443
rect 1066 6789 558846 7355
rect 1066 5701 558846 6267
rect 1066 4613 558846 5179
rect 1066 3525 558846 4091
rect 1066 2437 558846 3003
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 1104 8 559070 349840
<< metal2 >>
rect 3790 0 3846 800
rect 11058 0 11114 800
rect 18326 0 18382 800
rect 25594 0 25650 800
rect 32862 0 32918 800
rect 40130 0 40186 800
rect 47398 0 47454 800
rect 54666 0 54722 800
rect 61934 0 61990 800
rect 69202 0 69258 800
rect 76470 0 76526 800
rect 83738 0 83794 800
rect 91006 0 91062 800
rect 98274 0 98330 800
rect 105542 0 105598 800
rect 112810 0 112866 800
rect 120078 0 120134 800
rect 127346 0 127402 800
rect 134614 0 134670 800
rect 141882 0 141938 800
rect 149150 0 149206 800
rect 156418 0 156474 800
rect 163686 0 163742 800
rect 170954 0 171010 800
rect 178222 0 178278 800
rect 185490 0 185546 800
rect 192758 0 192814 800
rect 200026 0 200082 800
rect 207294 0 207350 800
rect 214562 0 214618 800
rect 221830 0 221886 800
rect 229098 0 229154 800
rect 236366 0 236422 800
rect 243634 0 243690 800
rect 250902 0 250958 800
rect 258170 0 258226 800
rect 265438 0 265494 800
rect 272706 0 272762 800
rect 279974 0 280030 800
rect 287242 0 287298 800
rect 294510 0 294566 800
rect 301778 0 301834 800
rect 309046 0 309102 800
rect 316314 0 316370 800
rect 323582 0 323638 800
rect 330850 0 330906 800
rect 338118 0 338174 800
rect 345386 0 345442 800
rect 352654 0 352710 800
rect 359922 0 359978 800
rect 367190 0 367246 800
rect 374458 0 374514 800
rect 381726 0 381782 800
rect 388994 0 389050 800
rect 396262 0 396318 800
rect 403530 0 403586 800
rect 410798 0 410854 800
rect 418066 0 418122 800
rect 425334 0 425390 800
rect 432602 0 432658 800
rect 439870 0 439926 800
rect 447138 0 447194 800
rect 454406 0 454462 800
rect 461674 0 461730 800
rect 468942 0 468998 800
rect 476210 0 476266 800
rect 483478 0 483534 800
rect 490746 0 490802 800
rect 498014 0 498070 800
rect 505282 0 505338 800
rect 512550 0 512606 800
rect 519818 0 519874 800
rect 527086 0 527142 800
rect 534354 0 534410 800
rect 541622 0 541678 800
rect 548890 0 548946 800
rect 556158 0 556214 800
<< obsm2 >>
rect 3792 856 559066 349829
rect 3902 2 11002 856
rect 11170 2 18270 856
rect 18438 2 25538 856
rect 25706 2 32806 856
rect 32974 2 40074 856
rect 40242 2 47342 856
rect 47510 2 54610 856
rect 54778 2 61878 856
rect 62046 2 69146 856
rect 69314 2 76414 856
rect 76582 2 83682 856
rect 83850 2 90950 856
rect 91118 2 98218 856
rect 98386 2 105486 856
rect 105654 2 112754 856
rect 112922 2 120022 856
rect 120190 2 127290 856
rect 127458 2 134558 856
rect 134726 2 141826 856
rect 141994 2 149094 856
rect 149262 2 156362 856
rect 156530 2 163630 856
rect 163798 2 170898 856
rect 171066 2 178166 856
rect 178334 2 185434 856
rect 185602 2 192702 856
rect 192870 2 199970 856
rect 200138 2 207238 856
rect 207406 2 214506 856
rect 214674 2 221774 856
rect 221942 2 229042 856
rect 229210 2 236310 856
rect 236478 2 243578 856
rect 243746 2 250846 856
rect 251014 2 258114 856
rect 258282 2 265382 856
rect 265550 2 272650 856
rect 272818 2 279918 856
rect 280086 2 287186 856
rect 287354 2 294454 856
rect 294622 2 301722 856
rect 301890 2 308990 856
rect 309158 2 316258 856
rect 316426 2 323526 856
rect 323694 2 330794 856
rect 330962 2 338062 856
rect 338230 2 345330 856
rect 345498 2 352598 856
rect 352766 2 359866 856
rect 360034 2 367134 856
rect 367302 2 374402 856
rect 374570 2 381670 856
rect 381838 2 388938 856
rect 389106 2 396206 856
rect 396374 2 403474 856
rect 403642 2 410742 856
rect 410910 2 418010 856
rect 418178 2 425278 856
rect 425446 2 432546 856
rect 432714 2 439814 856
rect 439982 2 447082 856
rect 447250 2 454350 856
rect 454518 2 461618 856
rect 461786 2 468886 856
rect 469054 2 476154 856
rect 476322 2 483422 856
rect 483590 2 490690 856
rect 490858 2 497958 856
rect 498126 2 505226 856
rect 505394 2 512494 856
rect 512662 2 519762 856
rect 519930 2 527030 856
rect 527198 2 534298 856
rect 534466 2 541566 856
rect 541734 2 548834 856
rect 549002 2 556102 856
rect 556270 2 559066 856
<< metal3 >>
rect 559200 344360 560000 344480
rect 559200 333480 560000 333600
rect 559200 322600 560000 322720
rect 559200 311720 560000 311840
rect 559200 300840 560000 300960
rect 559200 289960 560000 290080
rect 559200 279080 560000 279200
rect 559200 268200 560000 268320
rect 559200 257320 560000 257440
rect 559200 246440 560000 246560
rect 559200 235560 560000 235680
rect 559200 224680 560000 224800
rect 559200 213800 560000 213920
rect 559200 202920 560000 203040
rect 559200 192040 560000 192160
rect 559200 181160 560000 181280
rect 559200 170280 560000 170400
rect 559200 159400 560000 159520
rect 559200 148520 560000 148640
rect 559200 137640 560000 137760
rect 559200 126760 560000 126880
rect 559200 115880 560000 116000
rect 559200 105000 560000 105120
rect 559200 94120 560000 94240
rect 559200 83240 560000 83360
rect 559200 72360 560000 72480
rect 559200 61480 560000 61600
rect 559200 50600 560000 50720
rect 559200 39720 560000 39840
rect 559200 28840 560000 28960
rect 559200 17960 560000 18080
rect 559200 7080 560000 7200
<< obsm3 >>
rect 4210 344560 559200 349825
rect 4210 344280 559120 344560
rect 4210 333680 559200 344280
rect 4210 333400 559120 333680
rect 4210 322800 559200 333400
rect 4210 322520 559120 322800
rect 4210 311920 559200 322520
rect 4210 311640 559120 311920
rect 4210 301040 559200 311640
rect 4210 300760 559120 301040
rect 4210 290160 559200 300760
rect 4210 289880 559120 290160
rect 4210 279280 559200 289880
rect 4210 279000 559120 279280
rect 4210 268400 559200 279000
rect 4210 268120 559120 268400
rect 4210 257520 559200 268120
rect 4210 257240 559120 257520
rect 4210 246640 559200 257240
rect 4210 246360 559120 246640
rect 4210 235760 559200 246360
rect 4210 235480 559120 235760
rect 4210 224880 559200 235480
rect 4210 224600 559120 224880
rect 4210 214000 559200 224600
rect 4210 213720 559120 214000
rect 4210 203120 559200 213720
rect 4210 202840 559120 203120
rect 4210 192240 559200 202840
rect 4210 191960 559120 192240
rect 4210 181360 559200 191960
rect 4210 181080 559120 181360
rect 4210 170480 559200 181080
rect 4210 170200 559120 170480
rect 4210 159600 559200 170200
rect 4210 159320 559120 159600
rect 4210 148720 559200 159320
rect 4210 148440 559120 148720
rect 4210 137840 559200 148440
rect 4210 137560 559120 137840
rect 4210 126960 559200 137560
rect 4210 126680 559120 126960
rect 4210 116080 559200 126680
rect 4210 115800 559120 116080
rect 4210 105200 559200 115800
rect 4210 104920 559120 105200
rect 4210 94320 559200 104920
rect 4210 94040 559120 94320
rect 4210 83440 559200 94040
rect 4210 83160 559120 83440
rect 4210 72560 559200 83160
rect 4210 72280 559120 72560
rect 4210 61680 559200 72280
rect 4210 61400 559120 61680
rect 4210 50800 559200 61400
rect 4210 50520 559120 50800
rect 4210 39920 559200 50520
rect 4210 39640 559120 39920
rect 4210 29040 559200 39640
rect 4210 28760 559120 29040
rect 4210 18160 559200 28760
rect 4210 17880 559120 18160
rect 4210 7280 559200 17880
rect 4210 7000 559120 7280
rect 4210 35 559200 7000
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 139715 2048 142368 17101
rect 142848 2048 157728 17101
rect 158208 2048 173088 17101
rect 173568 2048 188448 17101
rect 188928 2048 203808 17101
rect 204288 2048 217061 17101
rect 139715 171 217061 2048
<< labels >>
rlabel metal2 s 250902 0 250958 800 6 irq[0]
port 1 nsew
rlabel metal2 s 258170 0 258226 800 6 irq[1]
port 2 nsew
rlabel metal2 s 265438 0 265494 800 6 irq[2]
port 3 nsew
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 4 nsew
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 4 nsew
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 4 nsew
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 4 nsew
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 4 nsew
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 4 nsew
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 4 nsew
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 4 nsew
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 4 nsew
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 4 nsew
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 4 nsew
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 4 nsew
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 4 nsew
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 4 nsew
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 4 nsew
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 4 nsew
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 4 nsew
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 4 nsew
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 4 nsew
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 5 nsew
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 5 nsew
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 5 nsew
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 5 nsew
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 5 nsew
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 5 nsew
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 5 nsew
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 5 nsew
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 5 nsew
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 5 nsew
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 5 nsew
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 5 nsew
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 5 nsew
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 5 nsew
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 5 nsew
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 5 nsew
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 5 nsew
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 5 nsew
rlabel metal2 s 3790 0 3846 800 6 wb_clk_i
port 6 nsew
rlabel metal2 s 11058 0 11114 800 6 wb_rst_i
port 7 nsew
rlabel metal2 s 323582 0 323638 800 6 wbs_ack_o
port 8 nsew
rlabel metal2 s 330850 0 330906 800 6 wbs_adr_i[0]
port 9 nsew
rlabel metal2 s 403530 0 403586 800 6 wbs_adr_i[10]
port 10 nsew
rlabel metal2 s 410798 0 410854 800 6 wbs_adr_i[11]
port 11 nsew
rlabel metal2 s 418066 0 418122 800 6 wbs_adr_i[12]
port 12 nsew
rlabel metal2 s 425334 0 425390 800 6 wbs_adr_i[13]
port 13 nsew
rlabel metal2 s 432602 0 432658 800 6 wbs_adr_i[14]
port 14 nsew
rlabel metal2 s 439870 0 439926 800 6 wbs_adr_i[15]
port 15 nsew
rlabel metal2 s 447138 0 447194 800 6 wbs_adr_i[16]
port 16 nsew
rlabel metal2 s 454406 0 454462 800 6 wbs_adr_i[17]
port 17 nsew
rlabel metal2 s 461674 0 461730 800 6 wbs_adr_i[18]
port 18 nsew
rlabel metal2 s 468942 0 468998 800 6 wbs_adr_i[19]
port 19 nsew
rlabel metal2 s 338118 0 338174 800 6 wbs_adr_i[1]
port 20 nsew
rlabel metal2 s 476210 0 476266 800 6 wbs_adr_i[20]
port 21 nsew
rlabel metal2 s 483478 0 483534 800 6 wbs_adr_i[21]
port 22 nsew
rlabel metal2 s 490746 0 490802 800 6 wbs_adr_i[22]
port 23 nsew
rlabel metal2 s 498014 0 498070 800 6 wbs_adr_i[23]
port 24 nsew
rlabel metal2 s 505282 0 505338 800 6 wbs_adr_i[24]
port 25 nsew
rlabel metal2 s 512550 0 512606 800 6 wbs_adr_i[25]
port 26 nsew
rlabel metal2 s 519818 0 519874 800 6 wbs_adr_i[26]
port 27 nsew
rlabel metal2 s 527086 0 527142 800 6 wbs_adr_i[27]
port 28 nsew
rlabel metal2 s 534354 0 534410 800 6 wbs_adr_i[28]
port 29 nsew
rlabel metal2 s 541622 0 541678 800 6 wbs_adr_i[29]
port 30 nsew
rlabel metal2 s 345386 0 345442 800 6 wbs_adr_i[2]
port 31 nsew
rlabel metal2 s 548890 0 548946 800 6 wbs_adr_i[30]
port 32 nsew
rlabel metal2 s 556158 0 556214 800 6 wbs_adr_i[31]
port 33 nsew
rlabel metal2 s 352654 0 352710 800 6 wbs_adr_i[3]
port 34 nsew
rlabel metal2 s 359922 0 359978 800 6 wbs_adr_i[4]
port 35 nsew
rlabel metal2 s 367190 0 367246 800 6 wbs_adr_i[5]
port 36 nsew
rlabel metal2 s 374458 0 374514 800 6 wbs_adr_i[6]
port 37 nsew
rlabel metal2 s 381726 0 381782 800 6 wbs_adr_i[7]
port 38 nsew
rlabel metal2 s 388994 0 389050 800 6 wbs_adr_i[8]
port 39 nsew
rlabel metal2 s 396262 0 396318 800 6 wbs_adr_i[9]
port 40 nsew
rlabel metal2 s 309046 0 309102 800 6 wbs_cyc_i
port 41 nsew
rlabel metal3 s 559200 7080 560000 7200 6 wbs_dat_i[0]
port 42 nsew
rlabel metal3 s 559200 115880 560000 116000 6 wbs_dat_i[10]
port 43 nsew
rlabel metal3 s 559200 126760 560000 126880 6 wbs_dat_i[11]
port 44 nsew
rlabel metal3 s 559200 137640 560000 137760 6 wbs_dat_i[12]
port 45 nsew
rlabel metal3 s 559200 148520 560000 148640 6 wbs_dat_i[13]
port 46 nsew
rlabel metal3 s 559200 159400 560000 159520 6 wbs_dat_i[14]
port 47 nsew
rlabel metal3 s 559200 170280 560000 170400 6 wbs_dat_i[15]
port 48 nsew
rlabel metal3 s 559200 181160 560000 181280 6 wbs_dat_i[16]
port 49 nsew
rlabel metal3 s 559200 192040 560000 192160 6 wbs_dat_i[17]
port 50 nsew
rlabel metal3 s 559200 202920 560000 203040 6 wbs_dat_i[18]
port 51 nsew
rlabel metal3 s 559200 213800 560000 213920 6 wbs_dat_i[19]
port 52 nsew
rlabel metal3 s 559200 17960 560000 18080 6 wbs_dat_i[1]
port 53 nsew
rlabel metal3 s 559200 224680 560000 224800 6 wbs_dat_i[20]
port 54 nsew
rlabel metal3 s 559200 235560 560000 235680 6 wbs_dat_i[21]
port 55 nsew
rlabel metal3 s 559200 246440 560000 246560 6 wbs_dat_i[22]
port 56 nsew
rlabel metal3 s 559200 257320 560000 257440 6 wbs_dat_i[23]
port 57 nsew
rlabel metal3 s 559200 268200 560000 268320 6 wbs_dat_i[24]
port 58 nsew
rlabel metal3 s 559200 279080 560000 279200 6 wbs_dat_i[25]
port 59 nsew
rlabel metal3 s 559200 289960 560000 290080 6 wbs_dat_i[26]
port 60 nsew
rlabel metal3 s 559200 300840 560000 300960 6 wbs_dat_i[27]
port 61 nsew
rlabel metal3 s 559200 311720 560000 311840 6 wbs_dat_i[28]
port 62 nsew
rlabel metal3 s 559200 322600 560000 322720 6 wbs_dat_i[29]
port 63 nsew
rlabel metal3 s 559200 28840 560000 28960 6 wbs_dat_i[2]
port 64 nsew
rlabel metal3 s 559200 333480 560000 333600 6 wbs_dat_i[30]
port 65 nsew
rlabel metal3 s 559200 344360 560000 344480 6 wbs_dat_i[31]
port 66 nsew
rlabel metal3 s 559200 39720 560000 39840 6 wbs_dat_i[3]
port 67 nsew
rlabel metal3 s 559200 50600 560000 50720 6 wbs_dat_i[4]
port 68 nsew
rlabel metal3 s 559200 61480 560000 61600 6 wbs_dat_i[5]
port 69 nsew
rlabel metal3 s 559200 72360 560000 72480 6 wbs_dat_i[6]
port 70 nsew
rlabel metal3 s 559200 83240 560000 83360 6 wbs_dat_i[7]
port 71 nsew
rlabel metal3 s 559200 94120 560000 94240 6 wbs_dat_i[8]
port 72 nsew
rlabel metal3 s 559200 105000 560000 105120 6 wbs_dat_i[9]
port 73 nsew
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[0]
port 74 nsew
rlabel metal2 s 91006 0 91062 800 6 wbs_dat_o[10]
port 75 nsew
rlabel metal2 s 98274 0 98330 800 6 wbs_dat_o[11]
port 76 nsew
rlabel metal2 s 105542 0 105598 800 6 wbs_dat_o[12]
port 77 nsew
rlabel metal2 s 112810 0 112866 800 6 wbs_dat_o[13]
port 78 nsew
rlabel metal2 s 120078 0 120134 800 6 wbs_dat_o[14]
port 79 nsew
rlabel metal2 s 127346 0 127402 800 6 wbs_dat_o[15]
port 80 nsew
rlabel metal2 s 134614 0 134670 800 6 wbs_dat_o[16]
port 81 nsew
rlabel metal2 s 141882 0 141938 800 6 wbs_dat_o[17]
port 82 nsew
rlabel metal2 s 149150 0 149206 800 6 wbs_dat_o[18]
port 83 nsew
rlabel metal2 s 156418 0 156474 800 6 wbs_dat_o[19]
port 84 nsew
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_o[1]
port 85 nsew
rlabel metal2 s 163686 0 163742 800 6 wbs_dat_o[20]
port 86 nsew
rlabel metal2 s 170954 0 171010 800 6 wbs_dat_o[21]
port 87 nsew
rlabel metal2 s 178222 0 178278 800 6 wbs_dat_o[22]
port 88 nsew
rlabel metal2 s 185490 0 185546 800 6 wbs_dat_o[23]
port 89 nsew
rlabel metal2 s 192758 0 192814 800 6 wbs_dat_o[24]
port 90 nsew
rlabel metal2 s 200026 0 200082 800 6 wbs_dat_o[25]
port 91 nsew
rlabel metal2 s 207294 0 207350 800 6 wbs_dat_o[26]
port 92 nsew
rlabel metal2 s 214562 0 214618 800 6 wbs_dat_o[27]
port 93 nsew
rlabel metal2 s 221830 0 221886 800 6 wbs_dat_o[28]
port 94 nsew
rlabel metal2 s 229098 0 229154 800 6 wbs_dat_o[29]
port 95 nsew
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[2]
port 96 nsew
rlabel metal2 s 236366 0 236422 800 6 wbs_dat_o[30]
port 97 nsew
rlabel metal2 s 243634 0 243690 800 6 wbs_dat_o[31]
port 98 nsew
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_o[3]
port 99 nsew
rlabel metal2 s 47398 0 47454 800 6 wbs_dat_o[4]
port 100 nsew
rlabel metal2 s 54666 0 54722 800 6 wbs_dat_o[5]
port 101 nsew
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_o[6]
port 102 nsew
rlabel metal2 s 69202 0 69258 800 6 wbs_dat_o[7]
port 103 nsew
rlabel metal2 s 76470 0 76526 800 6 wbs_dat_o[8]
port 104 nsew
rlabel metal2 s 83738 0 83794 800 6 wbs_dat_o[9]
port 105 nsew
rlabel metal2 s 272706 0 272762 800 6 wbs_sel_i[0]
port 106 nsew
rlabel metal2 s 279974 0 280030 800 6 wbs_sel_i[1]
port 107 nsew
rlabel metal2 s 287242 0 287298 800 6 wbs_sel_i[2]
port 108 nsew
rlabel metal2 s 294510 0 294566 800 6 wbs_sel_i[3]
port 109 nsew
rlabel metal2 s 301778 0 301834 800 6 wbs_stb_i
port 110 nsew
rlabel metal2 s 316314 0 316370 800 6 wbs_we_i
port 111 nsew
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 57010750
string GDS_FILE /home/nouran/user_proj_mul32/openlane/user_proj_mul32/runs/23_06_04_18_04/results/signoff/user_proj_mul32.magic.gds
string GDS_START 487258
<< end >>

