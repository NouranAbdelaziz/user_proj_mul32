magic
tech sky130B
magscale 1 2
timestamp 1676037725
use sky130_fd_pr__nfet_01v8__example_55959141808248  sky130_fd_pr__nfet_01v8__example_55959141808248_0
timestamp 1676037725
transform 1 0 910 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808445  sky130_fd_pr__nfet_01v8__example_55959141808445_0
timestamp 1676037725
transform 1 0 286 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_0
timestamp 1676037725
transform 1 0 442 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_1
timestamp 1676037725
transform 1 0 598 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_2
timestamp 1676037725
transform 1 0 754 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808455  sky130_fd_pr__nfet_01v8__example_55959141808455_0
timestamp 1676037725
transform -1 0 212 0 -1 1102
box -19 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808584  sky130_fd_pr__nfet_01v8__example_55959141808584_0
timestamp 1676037725
transform -1 0 212 0 -1 770
box 100 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808450  sky130_fd_pr__pfet_01v8__example_55959141808450_0
timestamp 1676037725
transform -1 0 720 0 -1 1650
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808451  sky130_fd_pr__pfet_01v8__example_55959141808451_0
timestamp 1676037725
transform 1 0 794 0 -1 1650
box -19 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808457  sky130_fd_pr__pfet_01v8__example_55959141808457_0
timestamp 1676037725
transform 1 0 72 0 -1 1650
box -1 0 297 1
<< properties >>
string GDS_END 43893042
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43878588
<< end >>
