magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< locali >>
rect 8981 8501 9015 8517
rect 8981 8451 9015 8467
rect 3290 7832 3324 7848
rect 3290 7782 3324 7798
rect 7517 7794 7551 7810
rect 7517 7744 7551 7760
rect 8981 7087 9015 7103
rect 6786 7053 8981 7087
rect 8981 7037 9015 7053
rect 3573 6790 3792 6824
rect 3758 6308 3792 6790
rect 5953 6380 5987 6396
rect 5953 6330 5987 6346
rect 3438 6191 3472 6207
rect 3438 6141 3472 6157
rect 3338 5943 3372 5959
rect 3338 5893 3372 5909
rect 8981 5673 9015 5689
rect 4504 5639 8981 5673
rect 8981 5623 9015 5639
rect 3305 5403 3339 5419
rect 3305 5353 3339 5369
rect 3438 5279 3472 5295
rect 3438 5229 3472 5245
rect 3571 5155 3605 5171
rect 3571 5105 3605 5121
rect 4101 4982 4135 4998
rect 4101 4932 4135 4948
rect 8981 4259 9015 4275
rect 4504 4225 8981 4259
rect 8981 4209 9015 4225
rect 4109 3536 4143 3552
rect 4109 3486 4143 3502
rect 3438 3363 3472 3379
rect 3438 3313 3472 3329
rect 3338 3115 3372 3131
rect 3338 3065 3372 3081
rect 8981 2845 9015 2861
rect 4620 2811 8981 2845
rect 8981 2795 9015 2811
rect 3555 2541 3740 2575
rect 3290 2176 3324 2192
rect 3555 2176 3589 2541
rect 3806 2327 3840 2343
rect 3806 2277 3840 2293
rect 3422 2142 3589 2176
rect 4477 2154 4511 2170
rect 3290 2126 3324 2142
rect 4477 2104 4511 2120
rect 8981 1431 9015 1447
rect 4988 1397 8981 1431
rect 8981 1381 9015 1397
rect 7299 724 7333 740
rect 3290 686 3324 702
rect 7299 674 7333 690
rect 3290 636 3324 652
rect 8981 17 9015 33
rect 8566 -17 8981 17
rect 8981 -33 9015 -17
<< viali >>
rect 8981 8467 9015 8501
rect 3290 7798 3324 7832
rect 7517 7760 7551 7794
rect 8981 7053 9015 7087
rect 5953 6346 5987 6380
rect 3438 6157 3472 6191
rect 3338 5909 3372 5943
rect 8981 5639 9015 5673
rect 3305 5369 3339 5403
rect 3438 5245 3472 5279
rect 3571 5121 3605 5155
rect 4101 4948 4135 4982
rect 8981 4225 9015 4259
rect 4109 3502 4143 3536
rect 3438 3329 3472 3363
rect 3338 3081 3372 3115
rect 8981 2811 9015 2845
rect 3806 2293 3840 2327
rect 3290 2142 3324 2176
rect 4477 2120 4511 2154
rect 8981 1397 9015 1431
rect 3290 652 3324 686
rect 7299 690 7333 724
rect 8981 -17 9015 17
<< metal1 >>
rect 8966 8458 8972 8510
rect 9024 8458 9030 8510
rect 2704 7789 2710 7841
rect 2762 7829 2768 7841
rect 3278 7832 3336 7838
rect 3278 7829 3290 7832
rect 2762 7801 3290 7829
rect 2762 7789 2768 7801
rect 3278 7798 3290 7801
rect 3324 7798 3336 7832
rect 3278 7792 3336 7798
rect 7502 7751 7508 7803
rect 7560 7751 7566 7803
rect 8966 7044 8972 7096
rect 9024 7044 9030 7096
rect 5938 6337 5944 6389
rect 5996 6337 6002 6389
rect 2620 6148 2626 6200
rect 2678 6188 2684 6200
rect 3426 6191 3484 6197
rect 3426 6188 3438 6191
rect 2678 6160 3438 6188
rect 2678 6148 2684 6160
rect 3426 6157 3438 6160
rect 3472 6157 3484 6191
rect 3426 6151 3484 6157
rect 2788 5900 2794 5952
rect 2846 5940 2852 5952
rect 3326 5943 3384 5949
rect 3326 5940 3338 5943
rect 2846 5912 3338 5940
rect 2846 5900 2852 5912
rect 3326 5909 3338 5912
rect 3372 5909 3384 5943
rect 3326 5903 3384 5909
rect 8966 5630 8972 5682
rect 9024 5630 9030 5682
rect 2620 5360 2626 5412
rect 2678 5400 2684 5412
rect 3293 5403 3351 5409
rect 3293 5400 3305 5403
rect 2678 5372 3305 5400
rect 2678 5360 2684 5372
rect 3293 5369 3305 5372
rect 3339 5369 3351 5403
rect 3293 5363 3351 5369
rect 2704 5236 2710 5288
rect 2762 5276 2768 5288
rect 3426 5279 3484 5285
rect 3426 5276 3438 5279
rect 2762 5248 3438 5276
rect 2762 5236 2768 5248
rect 3426 5245 3438 5248
rect 3472 5245 3484 5279
rect 3426 5239 3484 5245
rect 3040 5112 3046 5164
rect 3098 5152 3104 5164
rect 3559 5155 3617 5161
rect 3559 5152 3571 5155
rect 3098 5124 3571 5152
rect 3098 5112 3104 5124
rect 3559 5121 3571 5124
rect 3605 5121 3617 5155
rect 3559 5115 3617 5121
rect 4086 4939 4092 4991
rect 4144 4939 4150 4991
rect 1521 4296 1527 4348
rect 1579 4336 1585 4348
rect 2620 4336 2626 4348
rect 1579 4308 2626 4336
rect 1579 4296 1585 4308
rect 2620 4296 2626 4308
rect 2678 4296 2684 4348
rect 8966 4216 8972 4268
rect 9024 4216 9030 4268
rect 351 4136 357 4188
rect 409 4176 415 4188
rect 2872 4176 2878 4188
rect 409 4148 2878 4176
rect 409 4136 415 4148
rect 2872 4136 2878 4148
rect 2930 4136 2936 4188
rect 4094 3493 4100 3545
rect 4152 3493 4158 3545
rect 3040 3320 3046 3372
rect 3098 3360 3104 3372
rect 3426 3363 3484 3369
rect 3426 3360 3438 3363
rect 3098 3332 3438 3360
rect 3098 3320 3104 3332
rect 3426 3329 3438 3332
rect 3472 3329 3484 3363
rect 3426 3323 3484 3329
rect 2872 3072 2878 3124
rect 2930 3112 2936 3124
rect 3326 3115 3384 3121
rect 3326 3112 3338 3115
rect 2930 3084 3338 3112
rect 2930 3072 2936 3084
rect 3326 3081 3338 3084
rect 3372 3081 3384 3115
rect 3326 3075 3384 3081
rect 8966 2802 8972 2854
rect 9024 2802 9030 2854
rect 3791 2284 3797 2336
rect 3849 2284 3855 2336
rect 2872 2133 2878 2185
rect 2930 2173 2936 2185
rect 3278 2176 3336 2182
rect 3278 2173 3290 2176
rect 2930 2145 3290 2173
rect 2930 2133 2936 2145
rect 3278 2142 3290 2145
rect 3324 2142 3336 2176
rect 3278 2136 3336 2142
rect 4462 2111 4468 2163
rect 4520 2111 4526 2163
rect 8966 1388 8972 1440
rect 9024 1388 9030 1440
rect 3275 643 3281 695
rect 3333 643 3339 695
rect 7284 681 7290 733
rect 7342 681 7348 733
rect 8966 -26 8972 26
rect 9024 -26 9030 26
<< via1 >>
rect 8972 8501 9024 8510
rect 8972 8467 8981 8501
rect 8981 8467 9015 8501
rect 9015 8467 9024 8501
rect 8972 8458 9024 8467
rect 2710 7789 2762 7841
rect 7508 7794 7560 7803
rect 7508 7760 7517 7794
rect 7517 7760 7551 7794
rect 7551 7760 7560 7794
rect 7508 7751 7560 7760
rect 8972 7087 9024 7096
rect 8972 7053 8981 7087
rect 8981 7053 9015 7087
rect 9015 7053 9024 7087
rect 8972 7044 9024 7053
rect 5944 6380 5996 6389
rect 5944 6346 5953 6380
rect 5953 6346 5987 6380
rect 5987 6346 5996 6380
rect 5944 6337 5996 6346
rect 2626 6148 2678 6200
rect 2794 5900 2846 5952
rect 8972 5673 9024 5682
rect 8972 5639 8981 5673
rect 8981 5639 9015 5673
rect 9015 5639 9024 5673
rect 8972 5630 9024 5639
rect 2626 5360 2678 5412
rect 2710 5236 2762 5288
rect 3046 5112 3098 5164
rect 4092 4982 4144 4991
rect 4092 4948 4101 4982
rect 4101 4948 4135 4982
rect 4135 4948 4144 4982
rect 4092 4939 4144 4948
rect 1527 4296 1579 4348
rect 2626 4296 2678 4348
rect 8972 4259 9024 4268
rect 8972 4225 8981 4259
rect 8981 4225 9015 4259
rect 9015 4225 9024 4259
rect 8972 4216 9024 4225
rect 357 4136 409 4188
rect 2878 4136 2930 4188
rect 4100 3536 4152 3545
rect 4100 3502 4109 3536
rect 4109 3502 4143 3536
rect 4143 3502 4152 3536
rect 4100 3493 4152 3502
rect 3046 3320 3098 3372
rect 2878 3072 2930 3124
rect 8972 2845 9024 2854
rect 8972 2811 8981 2845
rect 8981 2811 9015 2845
rect 9015 2811 9024 2845
rect 8972 2802 9024 2811
rect 3797 2327 3849 2336
rect 3797 2293 3806 2327
rect 3806 2293 3840 2327
rect 3840 2293 3849 2327
rect 3797 2284 3849 2293
rect 2878 2133 2930 2185
rect 4468 2154 4520 2163
rect 4468 2120 4477 2154
rect 4477 2120 4511 2154
rect 4511 2120 4520 2154
rect 4468 2111 4520 2120
rect 8972 1431 9024 1440
rect 8972 1397 8981 1431
rect 8981 1397 9015 1431
rect 9015 1397 9024 1431
rect 8972 1388 9024 1397
rect 3281 686 3333 695
rect 3281 652 3290 686
rect 3290 652 3324 686
rect 3324 652 3333 686
rect 3281 643 3333 652
rect 7290 724 7342 733
rect 7290 690 7299 724
rect 7299 690 7333 724
rect 7333 690 7342 724
rect 7290 681 7342 690
rect 8972 17 9024 26
rect 8972 -17 8981 17
rect 8981 -17 9015 17
rect 9015 -17 9024 17
rect 8972 -26 9024 -17
<< metal2 >>
rect -57 17699 -29 17727
rect 1539 4354 1567 6401
rect 1527 4348 1579 4354
rect 1527 4290 1579 4296
rect 357 4188 409 4194
rect 357 4130 409 4136
rect 369 1414 397 4130
rect 1844 913 1900 922
rect 1844 848 1900 857
rect 137 538 203 590
rect 2350 531 2406 540
rect 2350 466 2406 475
rect 2554 0 2582 8524
rect 2638 6206 2666 8524
rect 2722 7847 2750 8524
rect 2710 7841 2762 7847
rect 2710 7783 2762 7789
rect 2626 6200 2678 6206
rect 2626 6142 2678 6148
rect 2638 5418 2666 6142
rect 2626 5412 2678 5418
rect 2626 5354 2678 5360
rect 2638 4354 2666 5354
rect 2722 5294 2750 7783
rect 2806 5958 2834 8524
rect 2794 5952 2846 5958
rect 2794 5894 2846 5900
rect 2710 5288 2762 5294
rect 2710 5230 2762 5236
rect 2626 4348 2678 4354
rect 2626 4290 2678 4296
rect 2638 0 2666 4290
rect 2722 1608 2750 5230
rect 2806 3556 2834 5894
rect 2890 4194 2918 8524
rect 2878 4188 2930 4194
rect 2878 4130 2930 4136
rect 2792 3547 2848 3556
rect 2792 3482 2848 3491
rect 2708 1599 2764 1608
rect 2708 1534 2764 1543
rect 2722 0 2750 1534
rect 2806 0 2834 3482
rect 2890 3130 2918 4130
rect 2878 3124 2930 3130
rect 2878 3066 2930 3072
rect 2890 2191 2918 3066
rect 2878 2185 2930 2191
rect 2878 2127 2930 2133
rect 2890 178 2918 2127
rect 2974 540 3002 8524
rect 3058 5170 3086 8524
rect 8970 8512 9026 8521
rect 8970 8447 9026 8456
rect 7508 7803 7560 7809
rect 7560 7763 9082 7791
rect 7508 7745 7560 7751
rect 8970 7098 9026 7107
rect 8970 7033 9026 7042
rect 5944 6389 5996 6395
rect 5996 6349 9082 6377
rect 5944 6331 5996 6337
rect 8970 5684 9026 5693
rect 8970 5619 9026 5628
rect 3046 5164 3098 5170
rect 3046 5106 3098 5112
rect 3058 3378 3086 5106
rect 4092 4991 4144 4997
rect 4144 4951 9082 4979
rect 4092 4933 4144 4939
rect 8970 4270 9026 4279
rect 8970 4205 9026 4214
rect 4098 3547 4154 3556
rect 4098 3482 4154 3491
rect 3046 3372 3098 3378
rect 3046 3314 3098 3320
rect 3058 2347 3086 3314
rect 8970 2856 9026 2865
rect 8970 2791 9026 2800
rect 3044 2338 3100 2347
rect 3044 2273 3100 2282
rect 3795 2338 3851 2347
rect 3795 2273 3851 2282
rect 3058 922 3086 2273
rect 4468 2163 4520 2169
rect 4468 2105 4520 2111
rect 4480 1608 4508 2105
rect 4466 1599 4522 1608
rect 4466 1534 4522 1543
rect 8970 1442 9026 1451
rect 8970 1377 9026 1386
rect 3044 913 3100 922
rect 3044 848 3100 857
rect 2960 531 3016 540
rect 2960 466 3016 475
rect 2876 169 2932 178
rect 2876 104 2932 113
rect 2890 0 2918 104
rect 2974 0 3002 466
rect 3058 0 3086 848
rect 7290 733 7342 739
rect 3281 695 3333 701
rect 7342 693 9082 721
rect 7290 675 7342 681
rect 3281 637 3333 643
rect 7302 178 7330 675
rect 7288 169 7344 178
rect 7288 104 7344 113
rect 8970 28 9026 37
rect 8970 -37 9026 -28
<< via2 >>
rect 1844 857 1900 913
rect 2350 475 2406 531
rect 2792 3491 2848 3547
rect 2708 1543 2764 1599
rect 8970 8510 9026 8512
rect 8970 8458 8972 8510
rect 8972 8458 9024 8510
rect 9024 8458 9026 8510
rect 8970 8456 9026 8458
rect 8970 7096 9026 7098
rect 8970 7044 8972 7096
rect 8972 7044 9024 7096
rect 9024 7044 9026 7096
rect 8970 7042 9026 7044
rect 8970 5682 9026 5684
rect 8970 5630 8972 5682
rect 8972 5630 9024 5682
rect 9024 5630 9026 5682
rect 8970 5628 9026 5630
rect 8970 4268 9026 4270
rect 8970 4216 8972 4268
rect 8972 4216 9024 4268
rect 9024 4216 9026 4268
rect 8970 4214 9026 4216
rect 4098 3545 4154 3547
rect 4098 3493 4100 3545
rect 4100 3493 4152 3545
rect 4152 3493 4154 3545
rect 4098 3491 4154 3493
rect 8970 2854 9026 2856
rect 8970 2802 8972 2854
rect 8972 2802 9024 2854
rect 9024 2802 9026 2854
rect 8970 2800 9026 2802
rect 3044 2282 3100 2338
rect 3795 2336 3851 2338
rect 3795 2284 3797 2336
rect 3797 2284 3849 2336
rect 3849 2284 3851 2336
rect 3795 2282 3851 2284
rect 4466 1543 4522 1599
rect 8970 1440 9026 1442
rect 8970 1388 8972 1440
rect 8972 1388 9024 1440
rect 9024 1388 9026 1440
rect 8970 1386 9026 1388
rect 3044 857 3100 913
rect 2960 475 3016 531
rect 2876 113 2932 169
rect 7288 113 7344 169
rect 8970 26 9026 28
rect 8970 -26 8972 26
rect 8972 -26 9024 26
rect 9024 -26 9026 26
rect 8970 -28 9026 -26
<< metal3 >>
rect 607 18333 705 18431
rect 1343 18333 1441 18431
rect 607 16919 705 17017
rect 1343 16919 1441 17017
rect 607 15505 705 15603
rect 1343 15505 1441 15603
rect 607 14091 705 14189
rect 1343 14091 1441 14189
rect 607 12677 705 12775
rect 1343 12677 1441 12775
rect 607 11263 705 11361
rect 1343 11263 1441 11361
rect 607 9849 705 9947
rect 1343 9849 1441 9947
rect 607 8435 705 8533
rect 1343 8435 1441 8533
rect 8949 8512 9047 8533
rect 8949 8456 8970 8512
rect 9026 8456 9047 8512
rect 8949 8435 9047 8456
rect 607 7021 705 7119
rect 1343 7021 1441 7119
rect 8949 7098 9047 7119
rect 8949 7042 8970 7098
rect 9026 7042 9047 7098
rect 8949 7021 9047 7042
rect 607 5607 705 5705
rect 1343 5607 1441 5705
rect 8949 5684 9047 5705
rect 8949 5628 8970 5684
rect 9026 5628 9047 5684
rect 8949 5607 9047 5628
rect 8949 4270 9047 4291
rect 8949 4214 8970 4270
rect 9026 4214 9047 4270
rect 8949 4193 9047 4214
rect 2787 3549 2853 3552
rect 4093 3549 4159 3552
rect 2787 3547 4159 3549
rect 2787 3491 2792 3547
rect 2848 3491 4098 3547
rect 4154 3491 4159 3547
rect 2787 3489 4159 3491
rect 2787 3486 2853 3489
rect 4093 3486 4159 3489
rect 8949 2856 9047 2877
rect 8949 2800 8970 2856
rect 9026 2800 9047 2856
rect 8949 2779 9047 2800
rect 3039 2340 3105 2343
rect 3790 2340 3856 2343
rect 3039 2338 3856 2340
rect 3039 2282 3044 2338
rect 3100 2282 3795 2338
rect 3851 2282 3856 2338
rect 3039 2280 3856 2282
rect 3039 2277 3105 2280
rect 3790 2277 3856 2280
rect 2703 1601 2769 1604
rect 4461 1601 4527 1604
rect 2703 1599 4527 1601
rect 2703 1543 2708 1599
rect 2764 1543 4466 1599
rect 4522 1543 4527 1599
rect 2703 1541 4527 1543
rect 2703 1538 2769 1541
rect 4461 1538 4527 1541
rect -49 1365 49 1463
rect 8949 1442 9047 1463
rect 8949 1386 8970 1442
rect 9026 1386 9047 1442
rect 8949 1365 9047 1386
rect 1839 915 1905 918
rect 3039 915 3105 918
rect 1839 913 3105 915
rect 1839 857 1844 913
rect 1900 857 3044 913
rect 3100 857 3105 913
rect 1839 855 3105 857
rect 1839 852 1905 855
rect 3039 852 3105 855
rect 2345 533 2411 536
rect 2955 533 3021 536
rect 2345 531 3021 533
rect 2345 475 2350 531
rect 2406 475 2960 531
rect 3016 475 3021 531
rect 2345 473 3021 475
rect 2345 470 2411 473
rect 2955 470 3021 473
rect 2871 171 2937 174
rect 7283 171 7349 174
rect 2871 169 7349 171
rect 2871 113 2876 169
rect 2932 113 7288 169
rect 7344 113 7349 169
rect 2871 111 7349 113
rect 2871 108 2937 111
rect 7283 108 7349 111
rect -49 -49 49 49
rect 8949 28 9047 49
rect 8949 -28 8970 28
rect 9026 -28 9047 28
rect 8949 -49 9047 -28
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_0
timestamp 1676037725
transform 1 0 8965 0 1 8447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_1
timestamp 1676037725
transform 1 0 8965 0 1 7033
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_2
timestamp 1676037725
transform 1 0 8965 0 1 5619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_3
timestamp 1676037725
transform 1 0 8965 0 1 7033
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_4
timestamp 1676037725
transform 1 0 8965 0 1 5619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_5
timestamp 1676037725
transform 1 0 8965 0 1 4205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_6
timestamp 1676037725
transform 1 0 8965 0 1 2791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_7
timestamp 1676037725
transform 1 0 8965 0 1 4205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_8
timestamp 1676037725
transform 1 0 8965 0 1 2791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_9
timestamp 1676037725
transform 1 0 8965 0 1 1377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_10
timestamp 1676037725
transform 1 0 8965 0 1 -37
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_11
timestamp 1676037725
transform 1 0 8965 0 1 1377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_12
timestamp 1676037725
transform 1 0 4093 0 1 3482
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_13
timestamp 1676037725
transform 1 0 3790 0 1 2273
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_14
timestamp 1676037725
transform 1 0 3790 0 1 2273
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_15
timestamp 1676037725
transform 1 0 2345 0 1 466
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_16
timestamp 1676037725
transform 1 0 1839 0 1 848
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_0
timestamp 1676037725
transform 1 0 8969 0 1 8451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1
timestamp 1676037725
transform 1 0 8969 0 1 7037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_2
timestamp 1676037725
transform 1 0 8969 0 1 5623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_3
timestamp 1676037725
transform 1 0 8969 0 1 7037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_4
timestamp 1676037725
transform 1 0 8969 0 1 5623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_5
timestamp 1676037725
transform 1 0 8969 0 1 4209
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_6
timestamp 1676037725
transform 1 0 8969 0 1 2795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_7
timestamp 1676037725
transform 1 0 8969 0 1 4209
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_8
timestamp 1676037725
transform 1 0 8969 0 1 2795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_9
timestamp 1676037725
transform 1 0 8969 0 1 1381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_10
timestamp 1676037725
transform 1 0 8969 0 1 -33
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_11
timestamp 1676037725
transform 1 0 8969 0 1 1381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_12
timestamp 1676037725
transform 1 0 5941 0 1 6330
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_13
timestamp 1676037725
transform 1 0 7505 0 1 7744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_14
timestamp 1676037725
transform 1 0 7287 0 1 674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_15
timestamp 1676037725
transform 1 0 7287 0 1 674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_16
timestamp 1676037725
transform 1 0 4097 0 1 3486
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_17
timestamp 1676037725
transform 1 0 4097 0 1 3486
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_18
timestamp 1676037725
transform 1 0 3426 0 1 3313
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_19
timestamp 1676037725
transform 1 0 3326 0 1 3065
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_20
timestamp 1676037725
transform 1 0 3794 0 1 2277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_21
timestamp 1676037725
transform 1 0 3794 0 1 2277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_22
timestamp 1676037725
transform 1 0 3278 0 1 2126
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_23
timestamp 1676037725
transform 1 0 3278 0 1 636
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_24
timestamp 1676037725
transform 1 0 3426 0 1 6141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_25
timestamp 1676037725
transform 1 0 3326 0 1 5893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_26
timestamp 1676037725
transform 1 0 4089 0 1 4932
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_27
timestamp 1676037725
transform 1 0 3559 0 1 5105
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_28
timestamp 1676037725
transform 1 0 3426 0 1 5229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_29
timestamp 1676037725
transform 1 0 3293 0 1 5353
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_30
timestamp 1676037725
transform 1 0 3278 0 1 7782
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_31
timestamp 1676037725
transform 1 0 4465 0 1 2104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1676037725
transform 1 0 8966 0 1 8452
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1676037725
transform 1 0 8966 0 1 7038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_2
timestamp 1676037725
transform 1 0 8966 0 1 5624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_3
timestamp 1676037725
transform 1 0 8966 0 1 7038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_4
timestamp 1676037725
transform 1 0 8966 0 1 5624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_5
timestamp 1676037725
transform 1 0 8966 0 1 4210
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_6
timestamp 1676037725
transform 1 0 8966 0 1 2796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_7
timestamp 1676037725
transform 1 0 8966 0 1 4210
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_8
timestamp 1676037725
transform 1 0 8966 0 1 2796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_9
timestamp 1676037725
transform 1 0 8966 0 1 1382
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_10
timestamp 1676037725
transform 1 0 8966 0 1 -32
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_11
timestamp 1676037725
transform 1 0 8966 0 1 1382
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_12
timestamp 1676037725
transform 1 0 7502 0 1 7745
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_13
timestamp 1676037725
transform 1 0 5938 0 1 6331
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_14
timestamp 1676037725
transform 1 0 7284 0 1 675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_15
timestamp 1676037725
transform 1 0 7284 0 1 675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_16
timestamp 1676037725
transform 1 0 4094 0 1 3487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_17
timestamp 1676037725
transform 1 0 4094 0 1 3487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_18
timestamp 1676037725
transform 1 0 3040 0 1 3314
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_19
timestamp 1676037725
transform 1 0 2872 0 1 3066
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_20
timestamp 1676037725
transform 1 0 3791 0 1 2278
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_21
timestamp 1676037725
transform 1 0 3791 0 1 2278
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_22
timestamp 1676037725
transform 1 0 2872 0 1 2127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_23
timestamp 1676037725
transform 1 0 3275 0 1 637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_24
timestamp 1676037725
transform 1 0 2620 0 1 6142
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_25
timestamp 1676037725
transform 1 0 2788 0 1 5894
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_26
timestamp 1676037725
transform 1 0 2620 0 1 4290
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_27
timestamp 1676037725
transform 1 0 1521 0 1 4290
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_28
timestamp 1676037725
transform 1 0 4086 0 1 4933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_29
timestamp 1676037725
transform 1 0 3040 0 1 5106
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_30
timestamp 1676037725
transform 1 0 2704 0 1 5230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_31
timestamp 1676037725
transform 1 0 2620 0 1 5354
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_32
timestamp 1676037725
transform 1 0 2704 0 1 7783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_33
timestamp 1676037725
transform 1 0 2872 0 1 4130
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_34
timestamp 1676037725
transform 1 0 351 0 1 4130
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_35
timestamp 1676037725
transform 1 0 4462 0 1 2105
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_0
timestamp 1676037725
transform 1 0 7283 0 1 104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_1
timestamp 1676037725
transform 1 0 2787 0 1 3482
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_2
timestamp 1676037725
transform 1 0 2703 0 1 1534
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_3
timestamp 1676037725
transform 1 0 3039 0 1 2273
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_4
timestamp 1676037725
transform 1 0 2871 0 1 104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_5
timestamp 1676037725
transform 1 0 2955 0 1 466
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_6
timestamp 1676037725
transform 1 0 3039 0 1 848
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_7
timestamp 1676037725
transform 1 0 4461 0 1 1534
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_delay_chain  sky130_sram_1kbyte_1rw1r_8x1024_8_delay_chain_0
timestamp 1676037725
transform 1 0 0 0 -1 18382
box -75 -49 1876 12783
use sky130_sram_1kbyte_1rw1r_8x1024_8_dff_buf_array_0  sky130_sram_1kbyte_1rw1r_8x1024_8_dff_buf_array_0_0
timestamp 1676037725
transform 1 0 0 0 1 0
box -49 -49 2590 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand2_0  sky130_sram_1kbyte_1rw1r_8x1024_8_pand2_0_0
timestamp 1676037725
transform 1 0 3226 0 1 2828
box -36 -17 1430 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand2_0  sky130_sram_1kbyte_1rw1r_8x1024_8_pand2_0_1
timestamp 1676037725
transform 1 0 3594 0 -1 2828
box -36 -17 1430 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_1  sky130_sram_1kbyte_1rw1r_8x1024_8_pand3_1_0
timestamp 1676037725
transform 1 0 3226 0 -1 5656
box -36 -17 1314 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_3  sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_3_0
timestamp 1676037725
transform 1 0 3226 0 -1 8484
box -36 -17 5808 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_6  sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_6_0
timestamp 1676037725
transform 1 0 3694 0 1 5656
box -36 -17 3128 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_7  sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_7_0
timestamp 1676037725
transform 1 0 3226 0 1 0
box -36 -17 5376 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_1  sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_1_0
timestamp 1676037725
transform 1 0 3226 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pnand2_1  sky130_sram_1kbyte_1rw1r_8x1024_8_pnand2_1_0
timestamp 1676037725
transform 1 0 3226 0 1 5656
box -36 -17 504 1471
<< labels >>
rlabel metal3 s -49 1365 49 1463 4 vdd
rlabel metal3 s 1343 5607 1441 5705 4 vdd
rlabel metal3 s 607 11263 705 11361 4 vdd
rlabel metal3 s 607 8435 705 8533 4 vdd
rlabel metal3 s 8949 7021 9047 7119 4 vdd
rlabel metal3 s 607 5607 705 5705 4 vdd
rlabel metal3 s 607 16919 705 17017 4 vdd
rlabel metal3 s 8949 4193 9047 4291 4 vdd
rlabel metal3 s 8949 1365 9047 1463 4 vdd
rlabel metal3 s 1343 16919 1441 17017 4 vdd
rlabel metal3 s 1343 8435 1441 8533 4 vdd
rlabel metal3 s 1343 11263 1441 11361 4 vdd
rlabel metal3 s 1343 14091 1441 14189 4 vdd
rlabel metal3 s 607 14091 705 14189 4 vdd
rlabel metal3 s 1343 9849 1441 9947 4 gnd
rlabel metal3 s 1343 15505 1441 15603 4 gnd
rlabel metal3 s 1343 12677 1441 12775 4 gnd
rlabel metal3 s 607 18333 705 18431 4 gnd
rlabel metal3 s 1343 18333 1441 18431 4 gnd
rlabel metal3 s 1343 7021 1441 7119 4 gnd
rlabel metal3 s 607 12677 705 12775 4 gnd
rlabel metal3 s 607 15505 705 15603 4 gnd
rlabel metal3 s 607 9849 705 9947 4 gnd
rlabel metal3 s -49 -49 49 49 4 gnd
rlabel metal3 s 8949 8435 9047 8533 4 gnd
rlabel metal3 s 607 7021 705 7119 4 gnd
rlabel metal3 s 8949 2779 9047 2877 4 gnd
rlabel metal3 s 8949 5607 9047 5705 4 gnd
rlabel metal3 s 8949 -49 9047 49 4 gnd
rlabel metal2 s 137 538 203 590 4 csb
rlabel metal2 s 7534 7763 9082 7791 4 wl_en
rlabel metal2 s 4118 4951 9082 4979 4 s_en
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
rlabel metal2 s 5970 6349 9082 6377 4 p_en_bar
rlabel metal2 s 3293 655 3321 683 4 clk
rlabel metal2 s 7316 693 9082 721 4 clk_buf
<< properties >>
string FIXED_BBOX 8965 -37 9031 0
string GDS_END 7083762
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 7063272
<< end >>
