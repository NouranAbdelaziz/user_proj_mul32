magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
rect 1478 5448 1524 5702
rect 2726 5448 2772 5702
rect 3974 5448 4020 5702
rect 5222 5448 5268 5702
rect 6470 5448 6516 5702
rect 7718 5448 7764 5702
rect 8966 5448 9012 5702
rect 10214 5448 10260 5702
rect 11462 5448 11508 5702
rect 12710 5448 12756 5702
rect 13958 5448 14004 5702
rect 15206 5448 15252 5702
rect 16454 5448 16500 5702
rect 17702 5448 17748 5702
rect 18950 5448 18996 5702
rect 20198 5448 20244 5702
rect 21446 5448 21492 5702
rect 22694 5448 22740 5702
rect 23942 5448 23988 5702
rect 25190 5448 25236 5702
rect 26438 5448 26484 5702
rect 27686 5448 27732 5702
rect 28934 5448 28980 5702
rect 30182 5448 30228 5702
rect 31430 5448 31476 5702
rect 32678 5448 32724 5702
rect 33926 5448 33972 5702
rect 35174 5448 35220 5702
rect 36422 5448 36468 5702
rect 37670 5448 37716 5702
rect 38918 5448 38964 5702
rect 40166 5448 40212 5702
rect 1573 3380 1601 3446
rect 1454 3352 1601 3380
rect 1454 2946 1482 3352
rect 1646 3300 1674 3446
rect 2821 3380 2849 3446
rect 2702 3352 2849 3380
rect 1646 3272 1946 3300
rect 1918 3070 1946 3272
rect 2702 2946 2730 3352
rect 2894 3300 2922 3446
rect 4069 3380 4097 3446
rect 3950 3352 4097 3380
rect 2894 3272 3194 3300
rect 3166 3070 3194 3272
rect 3950 2946 3978 3352
rect 4142 3300 4170 3446
rect 5317 3380 5345 3446
rect 5198 3352 5345 3380
rect 4142 3272 4442 3300
rect 4414 3070 4442 3272
rect 5198 2946 5226 3352
rect 5390 3300 5418 3446
rect 6565 3380 6593 3446
rect 6446 3352 6593 3380
rect 5390 3272 5690 3300
rect 5662 3070 5690 3272
rect 6446 2946 6474 3352
rect 6638 3300 6666 3446
rect 7813 3380 7841 3446
rect 7694 3352 7841 3380
rect 6638 3272 6938 3300
rect 6910 3070 6938 3272
rect 7694 2946 7722 3352
rect 7886 3300 7914 3446
rect 9061 3380 9089 3446
rect 8942 3352 9089 3380
rect 7886 3272 8186 3300
rect 8158 3070 8186 3272
rect 8942 2946 8970 3352
rect 9134 3300 9162 3446
rect 10309 3380 10337 3446
rect 10190 3352 10337 3380
rect 9134 3272 9434 3300
rect 9406 3070 9434 3272
rect 10190 2946 10218 3352
rect 10382 3300 10410 3446
rect 11557 3380 11585 3446
rect 11438 3352 11585 3380
rect 10382 3272 10682 3300
rect 10654 3070 10682 3272
rect 11438 2946 11466 3352
rect 11630 3300 11658 3446
rect 12805 3380 12833 3446
rect 12686 3352 12833 3380
rect 11630 3272 11930 3300
rect 11902 3070 11930 3272
rect 12686 2946 12714 3352
rect 12878 3300 12906 3446
rect 14053 3380 14081 3446
rect 13934 3352 14081 3380
rect 12878 3272 13178 3300
rect 13150 3070 13178 3272
rect 13934 2946 13962 3352
rect 14126 3300 14154 3446
rect 15301 3380 15329 3446
rect 15182 3352 15329 3380
rect 14126 3272 14426 3300
rect 14398 3070 14426 3272
rect 15182 2946 15210 3352
rect 15374 3300 15402 3446
rect 16549 3380 16577 3446
rect 16430 3352 16577 3380
rect 15374 3272 15674 3300
rect 15646 3070 15674 3272
rect 16430 2946 16458 3352
rect 16622 3300 16650 3446
rect 17797 3380 17825 3446
rect 17678 3352 17825 3380
rect 16622 3272 16922 3300
rect 16894 3070 16922 3272
rect 17678 2946 17706 3352
rect 17870 3300 17898 3446
rect 19045 3380 19073 3446
rect 18926 3352 19073 3380
rect 17870 3272 18170 3300
rect 18142 3070 18170 3272
rect 18926 2946 18954 3352
rect 19118 3300 19146 3446
rect 20293 3380 20321 3446
rect 20174 3352 20321 3380
rect 19118 3272 19418 3300
rect 19390 3070 19418 3272
rect 20174 2946 20202 3352
rect 20366 3300 20394 3446
rect 21541 3380 21569 3446
rect 21422 3352 21569 3380
rect 20366 3272 20666 3300
rect 20638 3070 20666 3272
rect 21422 2946 21450 3352
rect 21614 3300 21642 3446
rect 22789 3380 22817 3446
rect 22670 3352 22817 3380
rect 21614 3272 21914 3300
rect 21886 3070 21914 3272
rect 22670 2946 22698 3352
rect 22862 3300 22890 3446
rect 24037 3380 24065 3446
rect 23918 3352 24065 3380
rect 22862 3272 23162 3300
rect 23134 3070 23162 3272
rect 23918 2946 23946 3352
rect 24110 3300 24138 3446
rect 25285 3380 25313 3446
rect 25166 3352 25313 3380
rect 24110 3272 24410 3300
rect 24382 3070 24410 3272
rect 25166 2946 25194 3352
rect 25358 3300 25386 3446
rect 26533 3380 26561 3446
rect 26414 3352 26561 3380
rect 25358 3272 25658 3300
rect 25630 3070 25658 3272
rect 26414 2946 26442 3352
rect 26606 3300 26634 3446
rect 27781 3380 27809 3446
rect 27662 3352 27809 3380
rect 26606 3272 26906 3300
rect 26878 3070 26906 3272
rect 27662 2946 27690 3352
rect 27854 3300 27882 3446
rect 29029 3380 29057 3446
rect 28910 3352 29057 3380
rect 27854 3272 28154 3300
rect 28126 3070 28154 3272
rect 28910 2946 28938 3352
rect 29102 3300 29130 3446
rect 30277 3380 30305 3446
rect 30158 3352 30305 3380
rect 29102 3272 29402 3300
rect 29374 3070 29402 3272
rect 30158 2946 30186 3352
rect 30350 3300 30378 3446
rect 31525 3380 31553 3446
rect 31406 3352 31553 3380
rect 30350 3272 30650 3300
rect 30622 3070 30650 3272
rect 31406 2946 31434 3352
rect 31598 3300 31626 3446
rect 32773 3380 32801 3446
rect 32654 3352 32801 3380
rect 31598 3272 31898 3300
rect 31870 3070 31898 3272
rect 32654 2946 32682 3352
rect 32846 3300 32874 3446
rect 34021 3380 34049 3446
rect 33902 3352 34049 3380
rect 32846 3272 33146 3300
rect 33118 3070 33146 3272
rect 33902 2946 33930 3352
rect 34094 3300 34122 3446
rect 35269 3380 35297 3446
rect 35150 3352 35297 3380
rect 34094 3272 34394 3300
rect 34366 3070 34394 3272
rect 35150 2946 35178 3352
rect 35342 3300 35370 3446
rect 36517 3380 36545 3446
rect 36398 3352 36545 3380
rect 35342 3272 35642 3300
rect 35614 3070 35642 3272
rect 36398 2946 36426 3352
rect 36590 3300 36618 3446
rect 37765 3380 37793 3446
rect 37646 3352 37793 3380
rect 36590 3272 36890 3300
rect 36862 3070 36890 3272
rect 37646 2946 37674 3352
rect 37838 3300 37866 3446
rect 39013 3380 39041 3446
rect 38894 3352 39041 3380
rect 37838 3272 38138 3300
rect 38110 3070 38138 3272
rect 38894 2946 38922 3352
rect 39086 3300 39114 3446
rect 40261 3380 40289 3446
rect 40142 3352 40289 3380
rect 39086 3272 39386 3300
rect 39358 3070 39386 3272
rect 40142 2946 40170 3352
rect 40334 3300 40362 3446
rect 40334 3272 40634 3300
rect 40606 3070 40634 3272
rect 1454 1192 1482 1258
rect 1440 1164 1482 1192
rect 1440 252 1468 1164
rect 1918 1112 1946 1258
rect 1904 1084 1946 1112
rect 2050 1112 2078 1258
rect 2514 1192 2542 1258
rect 2702 1192 2730 1258
rect 2514 1164 2556 1192
rect 2050 1084 2092 1112
rect 1904 252 1932 1084
rect 2064 252 2092 1084
rect 2528 252 2556 1164
rect 2688 1164 2730 1192
rect 2688 252 2716 1164
rect 3166 1112 3194 1258
rect 3152 1084 3194 1112
rect 3298 1112 3326 1258
rect 3762 1192 3790 1258
rect 3950 1192 3978 1258
rect 3762 1164 3804 1192
rect 3298 1084 3340 1112
rect 3152 252 3180 1084
rect 3312 252 3340 1084
rect 3776 252 3804 1164
rect 3936 1164 3978 1192
rect 3936 252 3964 1164
rect 4414 1112 4442 1258
rect 4400 1084 4442 1112
rect 4546 1112 4574 1258
rect 5010 1192 5038 1258
rect 5198 1192 5226 1258
rect 5010 1164 5052 1192
rect 4546 1084 4588 1112
rect 4400 252 4428 1084
rect 4560 252 4588 1084
rect 5024 252 5052 1164
rect 5184 1164 5226 1192
rect 5184 252 5212 1164
rect 5662 1112 5690 1258
rect 5648 1084 5690 1112
rect 5794 1112 5822 1258
rect 6258 1192 6286 1258
rect 6446 1192 6474 1258
rect 6258 1164 6300 1192
rect 5794 1084 5836 1112
rect 5648 252 5676 1084
rect 5808 252 5836 1084
rect 6272 252 6300 1164
rect 6432 1164 6474 1192
rect 6432 252 6460 1164
rect 6910 1112 6938 1258
rect 6896 1084 6938 1112
rect 7042 1112 7070 1258
rect 7506 1192 7534 1258
rect 7694 1192 7722 1258
rect 7506 1164 7548 1192
rect 7042 1084 7084 1112
rect 6896 252 6924 1084
rect 7056 252 7084 1084
rect 7520 252 7548 1164
rect 7680 1164 7722 1192
rect 7680 252 7708 1164
rect 8158 1112 8186 1258
rect 8144 1084 8186 1112
rect 8290 1112 8318 1258
rect 8754 1192 8782 1258
rect 8942 1192 8970 1258
rect 8754 1164 8796 1192
rect 8290 1084 8332 1112
rect 8144 252 8172 1084
rect 8304 252 8332 1084
rect 8768 252 8796 1164
rect 8928 1164 8970 1192
rect 8928 252 8956 1164
rect 9406 1112 9434 1258
rect 9392 1084 9434 1112
rect 9538 1112 9566 1258
rect 10002 1192 10030 1258
rect 10190 1192 10218 1258
rect 10002 1164 10044 1192
rect 9538 1084 9580 1112
rect 9392 252 9420 1084
rect 9552 252 9580 1084
rect 10016 252 10044 1164
rect 10176 1164 10218 1192
rect 10176 252 10204 1164
rect 10654 1112 10682 1258
rect 10640 1084 10682 1112
rect 10786 1112 10814 1258
rect 11250 1192 11278 1258
rect 11438 1192 11466 1258
rect 11250 1164 11292 1192
rect 10786 1084 10828 1112
rect 10640 252 10668 1084
rect 10800 252 10828 1084
rect 11264 252 11292 1164
rect 11424 1164 11466 1192
rect 11424 252 11452 1164
rect 11902 1112 11930 1258
rect 11888 1084 11930 1112
rect 12034 1112 12062 1258
rect 12498 1192 12526 1258
rect 12686 1192 12714 1258
rect 12498 1164 12540 1192
rect 12034 1084 12076 1112
rect 11888 252 11916 1084
rect 12048 252 12076 1084
rect 12512 252 12540 1164
rect 12672 1164 12714 1192
rect 12672 252 12700 1164
rect 13150 1112 13178 1258
rect 13136 1084 13178 1112
rect 13282 1112 13310 1258
rect 13746 1192 13774 1258
rect 13934 1192 13962 1258
rect 13746 1164 13788 1192
rect 13282 1084 13324 1112
rect 13136 252 13164 1084
rect 13296 252 13324 1084
rect 13760 252 13788 1164
rect 13920 1164 13962 1192
rect 13920 252 13948 1164
rect 14398 1112 14426 1258
rect 14384 1084 14426 1112
rect 14530 1112 14558 1258
rect 14994 1192 15022 1258
rect 15182 1192 15210 1258
rect 14994 1164 15036 1192
rect 14530 1084 14572 1112
rect 14384 252 14412 1084
rect 14544 252 14572 1084
rect 15008 252 15036 1164
rect 15168 1164 15210 1192
rect 15168 252 15196 1164
rect 15646 1112 15674 1258
rect 15632 1084 15674 1112
rect 15778 1112 15806 1258
rect 16242 1192 16270 1258
rect 16430 1192 16458 1258
rect 16242 1164 16284 1192
rect 15778 1084 15820 1112
rect 15632 252 15660 1084
rect 15792 252 15820 1084
rect 16256 252 16284 1164
rect 16416 1164 16458 1192
rect 16416 252 16444 1164
rect 16894 1112 16922 1258
rect 16880 1084 16922 1112
rect 17026 1112 17054 1258
rect 17490 1192 17518 1258
rect 17678 1192 17706 1258
rect 17490 1164 17532 1192
rect 17026 1084 17068 1112
rect 16880 252 16908 1084
rect 17040 252 17068 1084
rect 17504 252 17532 1164
rect 17664 1164 17706 1192
rect 17664 252 17692 1164
rect 18142 1112 18170 1258
rect 18128 1084 18170 1112
rect 18274 1112 18302 1258
rect 18738 1192 18766 1258
rect 18926 1192 18954 1258
rect 18738 1164 18780 1192
rect 18274 1084 18316 1112
rect 18128 252 18156 1084
rect 18288 252 18316 1084
rect 18752 252 18780 1164
rect 18912 1164 18954 1192
rect 18912 252 18940 1164
rect 19390 1112 19418 1258
rect 19376 1084 19418 1112
rect 19522 1112 19550 1258
rect 19986 1192 20014 1258
rect 20174 1192 20202 1258
rect 19986 1164 20028 1192
rect 19522 1084 19564 1112
rect 19376 252 19404 1084
rect 19536 252 19564 1084
rect 20000 252 20028 1164
rect 20160 1164 20202 1192
rect 20160 252 20188 1164
rect 20638 1112 20666 1258
rect 20624 1084 20666 1112
rect 20770 1112 20798 1258
rect 21234 1192 21262 1258
rect 21422 1192 21450 1258
rect 21234 1164 21276 1192
rect 20770 1084 20812 1112
rect 20624 252 20652 1084
rect 20784 252 20812 1084
rect 21248 252 21276 1164
rect 21408 1164 21450 1192
rect 21408 252 21436 1164
rect 21886 1112 21914 1258
rect 21872 1084 21914 1112
rect 22018 1112 22046 1258
rect 22482 1192 22510 1258
rect 22670 1192 22698 1258
rect 22482 1164 22524 1192
rect 22018 1084 22060 1112
rect 21872 252 21900 1084
rect 22032 252 22060 1084
rect 22496 252 22524 1164
rect 22656 1164 22698 1192
rect 22656 252 22684 1164
rect 23134 1112 23162 1258
rect 23120 1084 23162 1112
rect 23266 1112 23294 1258
rect 23730 1192 23758 1258
rect 23918 1192 23946 1258
rect 23730 1164 23772 1192
rect 23266 1084 23308 1112
rect 23120 252 23148 1084
rect 23280 252 23308 1084
rect 23744 252 23772 1164
rect 23904 1164 23946 1192
rect 23904 252 23932 1164
rect 24382 1112 24410 1258
rect 24368 1084 24410 1112
rect 24514 1112 24542 1258
rect 24978 1192 25006 1258
rect 25166 1192 25194 1258
rect 24978 1164 25020 1192
rect 24514 1084 24556 1112
rect 24368 252 24396 1084
rect 24528 252 24556 1084
rect 24992 252 25020 1164
rect 25152 1164 25194 1192
rect 25152 252 25180 1164
rect 25630 1112 25658 1258
rect 25616 1084 25658 1112
rect 25762 1112 25790 1258
rect 26226 1192 26254 1258
rect 26414 1192 26442 1258
rect 26226 1164 26268 1192
rect 25762 1084 25804 1112
rect 25616 252 25644 1084
rect 25776 252 25804 1084
rect 26240 252 26268 1164
rect 26400 1164 26442 1192
rect 26400 252 26428 1164
rect 26878 1112 26906 1258
rect 26864 1084 26906 1112
rect 27010 1112 27038 1258
rect 27474 1192 27502 1258
rect 27662 1192 27690 1258
rect 27474 1164 27516 1192
rect 27010 1084 27052 1112
rect 26864 252 26892 1084
rect 27024 252 27052 1084
rect 27488 252 27516 1164
rect 27648 1164 27690 1192
rect 27648 252 27676 1164
rect 28126 1112 28154 1258
rect 28112 1084 28154 1112
rect 28258 1112 28286 1258
rect 28722 1192 28750 1258
rect 28910 1192 28938 1258
rect 28722 1164 28764 1192
rect 28258 1084 28300 1112
rect 28112 252 28140 1084
rect 28272 252 28300 1084
rect 28736 252 28764 1164
rect 28896 1164 28938 1192
rect 28896 252 28924 1164
rect 29374 1112 29402 1258
rect 29360 1084 29402 1112
rect 29506 1112 29534 1258
rect 29970 1192 29998 1258
rect 30158 1192 30186 1258
rect 29970 1164 30012 1192
rect 29506 1084 29548 1112
rect 29360 252 29388 1084
rect 29520 252 29548 1084
rect 29984 252 30012 1164
rect 30144 1164 30186 1192
rect 30144 252 30172 1164
rect 30622 1112 30650 1258
rect 30608 1084 30650 1112
rect 30754 1112 30782 1258
rect 31218 1192 31246 1258
rect 31406 1192 31434 1258
rect 31218 1164 31260 1192
rect 30754 1084 30796 1112
rect 30608 252 30636 1084
rect 30768 252 30796 1084
rect 31232 252 31260 1164
rect 31392 1164 31434 1192
rect 31392 252 31420 1164
rect 31870 1112 31898 1258
rect 31856 1084 31898 1112
rect 32002 1112 32030 1258
rect 32466 1192 32494 1258
rect 32654 1192 32682 1258
rect 32466 1164 32508 1192
rect 32002 1084 32044 1112
rect 31856 252 31884 1084
rect 32016 252 32044 1084
rect 32480 252 32508 1164
rect 32640 1164 32682 1192
rect 32640 252 32668 1164
rect 33118 1112 33146 1258
rect 33104 1084 33146 1112
rect 33250 1112 33278 1258
rect 33714 1192 33742 1258
rect 33902 1192 33930 1258
rect 33714 1164 33756 1192
rect 33250 1084 33292 1112
rect 33104 252 33132 1084
rect 33264 252 33292 1084
rect 33728 252 33756 1164
rect 33888 1164 33930 1192
rect 33888 252 33916 1164
rect 34366 1112 34394 1258
rect 34352 1084 34394 1112
rect 34498 1112 34526 1258
rect 34962 1192 34990 1258
rect 35150 1192 35178 1258
rect 34962 1164 35004 1192
rect 34498 1084 34540 1112
rect 34352 252 34380 1084
rect 34512 252 34540 1084
rect 34976 252 35004 1164
rect 35136 1164 35178 1192
rect 35136 252 35164 1164
rect 35614 1112 35642 1258
rect 35600 1084 35642 1112
rect 35746 1112 35774 1258
rect 36210 1192 36238 1258
rect 36398 1192 36426 1258
rect 36210 1164 36252 1192
rect 35746 1084 35788 1112
rect 35600 252 35628 1084
rect 35760 252 35788 1084
rect 36224 252 36252 1164
rect 36384 1164 36426 1192
rect 36384 252 36412 1164
rect 36862 1112 36890 1258
rect 36848 1084 36890 1112
rect 36994 1112 37022 1258
rect 37458 1192 37486 1258
rect 37646 1192 37674 1258
rect 37458 1164 37500 1192
rect 36994 1084 37036 1112
rect 36848 252 36876 1084
rect 37008 252 37036 1084
rect 37472 252 37500 1164
rect 37632 1164 37674 1192
rect 37632 252 37660 1164
rect 38110 1112 38138 1258
rect 38096 1084 38138 1112
rect 38242 1112 38270 1258
rect 38706 1192 38734 1258
rect 38894 1192 38922 1258
rect 38706 1164 38748 1192
rect 38242 1084 38284 1112
rect 38096 252 38124 1084
rect 38256 252 38284 1084
rect 38720 252 38748 1164
rect 38880 1164 38922 1192
rect 38880 252 38908 1164
rect 39358 1112 39386 1258
rect 39344 1084 39386 1112
rect 39490 1112 39518 1258
rect 39954 1192 39982 1258
rect 40142 1192 40170 1258
rect 39954 1164 39996 1192
rect 39490 1084 39532 1112
rect 39344 252 39372 1084
rect 39504 252 39532 1084
rect 39968 252 39996 1164
rect 40128 1164 40170 1192
rect 40128 252 40156 1164
rect 40606 1112 40634 1258
rect 40592 1084 40634 1112
rect 40738 1112 40766 1258
rect 41202 1192 41230 1258
rect 41202 1164 41244 1192
rect 40738 1084 40780 1112
rect 40592 252 40620 1084
rect 40752 252 40780 1084
rect 41216 252 41244 1164
rect 41376 252 41404 1006
rect 41840 252 41868 1006
<< metal3 >>
rect 1706 5545 1804 5643
rect 2954 5545 3052 5643
rect 4202 5545 4300 5643
rect 5450 5545 5548 5643
rect 6698 5545 6796 5643
rect 7946 5545 8044 5643
rect 9194 5545 9292 5643
rect 10442 5545 10540 5643
rect 11690 5545 11788 5643
rect 12938 5545 13036 5643
rect 14186 5545 14284 5643
rect 15434 5545 15532 5643
rect 16682 5545 16780 5643
rect 17930 5545 18028 5643
rect 19178 5545 19276 5643
rect 20426 5545 20524 5643
rect 21674 5545 21772 5643
rect 22922 5545 23020 5643
rect 24170 5545 24268 5643
rect 25418 5545 25516 5643
rect 26666 5545 26764 5643
rect 27914 5545 28012 5643
rect 29162 5545 29260 5643
rect 30410 5545 30508 5643
rect 31658 5545 31756 5643
rect 32906 5545 33004 5643
rect 34154 5545 34252 5643
rect 35402 5545 35500 5643
rect 36650 5545 36748 5643
rect 37898 5545 37996 5643
rect 39146 5545 39244 5643
rect 40394 5545 40492 5643
rect 1706 5223 1804 5321
rect 2954 5223 3052 5321
rect 4202 5223 4300 5321
rect 5450 5223 5548 5321
rect 6698 5223 6796 5321
rect 7946 5223 8044 5321
rect 9194 5223 9292 5321
rect 10442 5223 10540 5321
rect 11690 5223 11788 5321
rect 12938 5223 13036 5321
rect 14186 5223 14284 5321
rect 15434 5223 15532 5321
rect 16682 5223 16780 5321
rect 17930 5223 18028 5321
rect 19178 5223 19276 5321
rect 20426 5223 20524 5321
rect 21674 5223 21772 5321
rect 22922 5223 23020 5321
rect 24170 5223 24268 5321
rect 25418 5223 25516 5321
rect 26666 5223 26764 5321
rect 27914 5223 28012 5321
rect 29162 5223 29260 5321
rect 30410 5223 30508 5321
rect 31658 5223 31756 5321
rect 32906 5223 33004 5321
rect 34154 5223 34252 5321
rect 35402 5223 35500 5321
rect 36650 5223 36748 5321
rect 37898 5223 37996 5321
rect 39146 5223 39244 5321
rect 40394 5223 40492 5321
rect 1694 4385 1792 4483
rect 2942 4385 3040 4483
rect 4190 4385 4288 4483
rect 5438 4385 5536 4483
rect 6686 4385 6784 4483
rect 7934 4385 8032 4483
rect 9182 4385 9280 4483
rect 10430 4385 10528 4483
rect 11678 4385 11776 4483
rect 12926 4385 13024 4483
rect 14174 4385 14272 4483
rect 15422 4385 15520 4483
rect 16670 4385 16768 4483
rect 17918 4385 18016 4483
rect 19166 4385 19264 4483
rect 20414 4385 20512 4483
rect 21662 4385 21760 4483
rect 22910 4385 23008 4483
rect 24158 4385 24256 4483
rect 25406 4385 25504 4483
rect 26654 4385 26752 4483
rect 27902 4385 28000 4483
rect 29150 4385 29248 4483
rect 30398 4385 30496 4483
rect 31646 4385 31744 4483
rect 32894 4385 32992 4483
rect 34142 4385 34240 4483
rect 35390 4385 35488 4483
rect 36638 4385 36736 4483
rect 37886 4385 37984 4483
rect 39134 4385 39232 4483
rect 40382 4385 40480 4483
rect 1776 3611 1874 3709
rect 3024 3611 3122 3709
rect 4272 3611 4370 3709
rect 5520 3611 5618 3709
rect 6768 3611 6866 3709
rect 8016 3611 8114 3709
rect 9264 3611 9362 3709
rect 10512 3611 10610 3709
rect 11760 3611 11858 3709
rect 13008 3611 13106 3709
rect 14256 3611 14354 3709
rect 15504 3611 15602 3709
rect 16752 3611 16850 3709
rect 18000 3611 18098 3709
rect 19248 3611 19346 3709
rect 20496 3611 20594 3709
rect 21744 3611 21842 3709
rect 22992 3611 23090 3709
rect 24240 3611 24338 3709
rect 25488 3611 25586 3709
rect 26736 3611 26834 3709
rect 27984 3611 28082 3709
rect 29232 3611 29330 3709
rect 30480 3611 30578 3709
rect 31728 3611 31826 3709
rect 32976 3611 33074 3709
rect 34224 3611 34322 3709
rect 35472 3611 35570 3709
rect 36720 3611 36818 3709
rect 37968 3611 38066 3709
rect 39216 3611 39314 3709
rect 40464 3611 40562 3709
rect 0 3478 40562 3538
rect 0 2762 41310 2822
rect 0 2638 41310 2698
rect 1949 1862 2047 1960
rect 3197 1862 3295 1960
rect 4445 1862 4543 1960
rect 5693 1862 5791 1960
rect 6941 1862 7039 1960
rect 8189 1862 8287 1960
rect 9437 1862 9535 1960
rect 10685 1862 10783 1960
rect 11933 1862 12031 1960
rect 13181 1862 13279 1960
rect 14429 1862 14527 1960
rect 15677 1862 15775 1960
rect 16925 1862 17023 1960
rect 18173 1862 18271 1960
rect 19421 1862 19519 1960
rect 20669 1862 20767 1960
rect 21917 1862 22015 1960
rect 23165 1862 23263 1960
rect 24413 1862 24511 1960
rect 25661 1862 25759 1960
rect 26909 1862 27007 1960
rect 28157 1862 28255 1960
rect 29405 1862 29503 1960
rect 30653 1862 30751 1960
rect 31901 1862 31999 1960
rect 33149 1862 33247 1960
rect 34397 1862 34495 1960
rect 35645 1862 35743 1960
rect 36893 1862 36991 1960
rect 38141 1862 38239 1960
rect 39389 1862 39487 1960
rect 40637 1862 40735 1960
rect 0 951 41934 1011
rect 1518 313 1616 411
rect 2380 313 2478 411
rect 2766 313 2864 411
rect 3628 313 3726 411
rect 4014 313 4112 411
rect 4876 313 4974 411
rect 5262 313 5360 411
rect 6124 313 6222 411
rect 6510 313 6608 411
rect 7372 313 7470 411
rect 7758 313 7856 411
rect 8620 313 8718 411
rect 9006 313 9104 411
rect 9868 313 9966 411
rect 10254 313 10352 411
rect 11116 313 11214 411
rect 11502 313 11600 411
rect 12364 313 12462 411
rect 12750 313 12848 411
rect 13612 313 13710 411
rect 13998 313 14096 411
rect 14860 313 14958 411
rect 15246 313 15344 411
rect 16108 313 16206 411
rect 16494 313 16592 411
rect 17356 313 17454 411
rect 17742 313 17840 411
rect 18604 313 18702 411
rect 18990 313 19088 411
rect 19852 313 19950 411
rect 20238 313 20336 411
rect 21100 313 21198 411
rect 21486 313 21584 411
rect 22348 313 22446 411
rect 22734 313 22832 411
rect 23596 313 23694 411
rect 23982 313 24080 411
rect 24844 313 24942 411
rect 25230 313 25328 411
rect 26092 313 26190 411
rect 26478 313 26576 411
rect 27340 313 27438 411
rect 27726 313 27824 411
rect 28588 313 28686 411
rect 28974 313 29072 411
rect 29836 313 29934 411
rect 30222 313 30320 411
rect 31084 313 31182 411
rect 31470 313 31568 411
rect 32332 313 32430 411
rect 32718 313 32816 411
rect 33580 313 33678 411
rect 33966 313 34064 411
rect 34828 313 34926 411
rect 35214 313 35312 411
rect 36076 313 36174 411
rect 36462 313 36560 411
rect 37324 313 37422 411
rect 37710 313 37808 411
rect 38572 313 38670 411
rect 38958 313 39056 411
rect 39820 313 39918 411
rect 40206 313 40304 411
rect 41068 313 41166 411
rect 41454 313 41552 411
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array_0  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array_0_0
timestamp 1676037725
transform 1 0 0 0 -1 3194
box 0 87 41310 1936
use sky130_sram_1kbyte_1rw1r_32x256_8_precharge_array_0  sky130_sram_1kbyte_1rw1r_32x256_8_precharge_array_0_0
timestamp 1676037725
transform 1 0 0 0 -1 1006
box 0 -12 41934 768
use sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array  sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0
timestamp 1676037725
transform 1 0 0 0 -1 5702
box 0 0 40999 2256
<< labels >>
rlabel metal3 s 26654 4385 26752 4483 4 vdd
rlabel metal3 s 22922 5223 23020 5321 4 vdd
rlabel metal3 s 25418 5223 25516 5321 4 vdd
rlabel metal3 s 40394 5223 40492 5321 4 vdd
rlabel metal3 s 30410 5223 30508 5321 4 vdd
rlabel metal3 s 37886 4385 37984 4483 4 vdd
rlabel metal3 s 22910 4385 23008 4483 4 vdd
rlabel metal3 s 26666 5223 26764 5321 4 vdd
rlabel metal3 s 32894 4385 32992 4483 4 vdd
rlabel metal3 s 37898 5223 37996 5321 4 vdd
rlabel metal3 s 32906 5223 33004 5321 4 vdd
rlabel metal3 s 27914 5223 28012 5321 4 vdd
rlabel metal3 s 35390 4385 35488 4483 4 vdd
rlabel metal3 s 21674 5223 21772 5321 4 vdd
rlabel metal3 s 29150 4385 29248 4483 4 vdd
rlabel metal3 s 34142 4385 34240 4483 4 vdd
rlabel metal3 s 27902 4385 28000 4483 4 vdd
rlabel metal3 s 39146 5223 39244 5321 4 vdd
rlabel metal3 s 25406 4385 25504 4483 4 vdd
rlabel metal3 s 36650 5223 36748 5321 4 vdd
rlabel metal3 s 31646 4385 31744 4483 4 vdd
rlabel metal3 s 29162 5223 29260 5321 4 vdd
rlabel metal3 s 31658 5223 31756 5321 4 vdd
rlabel metal3 s 21662 4385 21760 4483 4 vdd
rlabel metal3 s 24170 5223 24268 5321 4 vdd
rlabel metal3 s 40382 4385 40480 4483 4 vdd
rlabel metal3 s 36638 4385 36736 4483 4 vdd
rlabel metal3 s 30398 4385 30496 4483 4 vdd
rlabel metal3 s 34154 5223 34252 5321 4 vdd
rlabel metal3 s 35402 5223 35500 5321 4 vdd
rlabel metal3 s 39134 4385 39232 4483 4 vdd
rlabel metal3 s 24158 4385 24256 4483 4 vdd
rlabel metal3 s 34224 3611 34322 3709 4 gnd
rlabel metal3 s 30410 5545 30508 5643 4 gnd
rlabel metal3 s 34397 1862 34495 1960 4 gnd
rlabel metal3 s 39146 5545 39244 5643 4 gnd
rlabel metal3 s 26736 3611 26834 3709 4 gnd
rlabel metal3 s 35402 5545 35500 5643 4 gnd
rlabel metal3 s 22922 5545 23020 5643 4 gnd
rlabel metal3 s 29162 5545 29260 5643 4 gnd
rlabel metal3 s 36720 3611 36818 3709 4 gnd
rlabel metal3 s 31728 3611 31826 3709 4 gnd
rlabel metal3 s 36650 5545 36748 5643 4 gnd
rlabel metal3 s 24170 5545 24268 5643 4 gnd
rlabel metal3 s 21917 1862 22015 1960 4 gnd
rlabel metal3 s 21744 3611 21842 3709 4 gnd
rlabel metal3 s 27914 5545 28012 5643 4 gnd
rlabel metal3 s 23165 1862 23263 1960 4 gnd
rlabel metal3 s 40637 1862 40735 1960 4 gnd
rlabel metal3 s 22992 3611 23090 3709 4 gnd
rlabel metal3 s 21674 5545 21772 5643 4 gnd
rlabel metal3 s 29405 1862 29503 1960 4 gnd
rlabel metal3 s 33149 1862 33247 1960 4 gnd
rlabel metal3 s 25418 5545 25516 5643 4 gnd
rlabel metal3 s 34154 5545 34252 5643 4 gnd
rlabel metal3 s 24413 1862 24511 1960 4 gnd
rlabel metal3 s 26666 5545 26764 5643 4 gnd
rlabel metal3 s 24240 3611 24338 3709 4 gnd
rlabel metal3 s 25661 1862 25759 1960 4 gnd
rlabel metal3 s 36893 1862 36991 1960 4 gnd
rlabel metal3 s 38141 1862 38239 1960 4 gnd
rlabel metal3 s 40464 3611 40562 3709 4 gnd
rlabel metal3 s 37898 5545 37996 5643 4 gnd
rlabel metal3 s 25488 3611 25586 3709 4 gnd
rlabel metal3 s 26909 1862 27007 1960 4 gnd
rlabel metal3 s 35645 1862 35743 1960 4 gnd
rlabel metal3 s 31901 1862 31999 1960 4 gnd
rlabel metal3 s 31658 5545 31756 5643 4 gnd
rlabel metal3 s 32976 3611 33074 3709 4 gnd
rlabel metal3 s 32906 5545 33004 5643 4 gnd
rlabel metal3 s 29232 3611 29330 3709 4 gnd
rlabel metal3 s 30653 1862 30751 1960 4 gnd
rlabel metal3 s 28157 1862 28255 1960 4 gnd
rlabel metal3 s 39389 1862 39487 1960 4 gnd
rlabel metal3 s 37968 3611 38066 3709 4 gnd
rlabel metal3 s 30480 3611 30578 3709 4 gnd
rlabel metal3 s 27984 3611 28082 3709 4 gnd
rlabel metal3 s 39216 3611 39314 3709 4 gnd
rlabel metal3 s 35472 3611 35570 3709 4 gnd
rlabel metal3 s 40394 5545 40492 5643 4 gnd
rlabel metal3 s 19248 3611 19346 3709 4 gnd
rlabel metal3 s 16670 4385 16768 4483 4 vdd
rlabel metal3 s 14186 5545 14284 5643 4 gnd
rlabel metal3 s 1694 4385 1792 4483 4 vdd
rlabel metal3 s 6698 5223 6796 5321 4 vdd
rlabel metal3 s 18000 3611 18098 3709 4 gnd
rlabel metal3 s 9264 3611 9362 3709 4 gnd
rlabel metal3 s 4202 5223 4300 5321 4 vdd
rlabel metal3 s 20414 4385 20512 4483 4 vdd
rlabel metal3 s 9194 5223 9292 5321 4 vdd
rlabel metal3 s 16752 3611 16850 3709 4 gnd
rlabel metal3 s 19166 4385 19264 4483 4 vdd
rlabel metal3 s 5520 3611 5618 3709 4 gnd
rlabel metal3 s 10430 4385 10528 4483 4 vdd
rlabel metal3 s 15422 4385 15520 4483 4 vdd
rlabel metal3 s 7934 4385 8032 4483 4 vdd
rlabel metal3 s 0 3478 40562 3538 4 s_en
rlabel metal3 s 19421 1862 19519 1960 4 gnd
rlabel metal3 s 8189 1862 8287 1960 4 gnd
rlabel metal3 s 19178 5223 19276 5321 4 vdd
rlabel metal3 s 6768 3611 6866 3709 4 gnd
rlabel metal3 s 17930 5223 18028 5321 4 vdd
rlabel metal3 s 16682 5223 16780 5321 4 vdd
rlabel metal3 s 2954 5223 3052 5321 4 vdd
rlabel metal3 s 12926 4385 13024 4483 4 vdd
rlabel metal3 s 12938 5223 13036 5321 4 vdd
rlabel metal3 s 11690 5545 11788 5643 4 gnd
rlabel metal3 s 0 951 41934 1011 4 p_en_bar
rlabel metal3 s 4202 5545 4300 5643 4 gnd
rlabel metal3 s 11933 1862 12031 1960 4 gnd
rlabel metal3 s 17918 4385 18016 4483 4 vdd
rlabel metal3 s 10442 5223 10540 5321 4 vdd
rlabel metal3 s 7946 5545 8044 5643 4 gnd
rlabel metal3 s 6686 4385 6784 4483 4 vdd
rlabel metal3 s 20669 1862 20767 1960 4 gnd
rlabel metal3 s 14256 3611 14354 3709 4 gnd
rlabel metal3 s 7946 5223 8044 5321 4 vdd
rlabel metal3 s 18173 1862 18271 1960 4 gnd
rlabel metal3 s 15434 5223 15532 5321 4 vdd
rlabel metal3 s 2942 4385 3040 4483 4 vdd
rlabel metal3 s 20426 5223 20524 5321 4 vdd
rlabel metal3 s 10442 5545 10540 5643 4 gnd
rlabel metal3 s 14429 1862 14527 1960 4 gnd
rlabel metal3 s 12938 5545 13036 5643 4 gnd
rlabel metal3 s 4190 4385 4288 4483 4 vdd
rlabel metal3 s 14186 5223 14284 5321 4 vdd
rlabel metal3 s 6941 1862 7039 1960 4 gnd
rlabel metal3 s 10685 1862 10783 1960 4 gnd
rlabel metal3 s 4445 1862 4543 1960 4 gnd
rlabel metal3 s 1949 1862 2047 1960 4 gnd
rlabel metal3 s 5438 4385 5536 4483 4 vdd
rlabel metal3 s 1706 5223 1804 5321 4 vdd
rlabel metal3 s 16925 1862 17023 1960 4 gnd
rlabel metal3 s 11678 4385 11776 4483 4 vdd
rlabel metal3 s 5450 5223 5548 5321 4 vdd
rlabel metal3 s 4272 3611 4370 3709 4 gnd
rlabel metal3 s 19178 5545 19276 5643 4 gnd
rlabel metal3 s 11690 5223 11788 5321 4 vdd
rlabel metal3 s 5693 1862 5791 1960 4 gnd
rlabel metal3 s 0 2762 41310 2822 4 sel_0
rlabel metal3 s 15504 3611 15602 3709 4 gnd
rlabel metal3 s 0 2638 41310 2698 4 sel_1
rlabel metal3 s 1776 3611 1874 3709 4 gnd
rlabel metal3 s 20496 3611 20594 3709 4 gnd
rlabel metal3 s 9437 1862 9535 1960 4 gnd
rlabel metal3 s 1706 5545 1804 5643 4 gnd
rlabel metal3 s 13181 1862 13279 1960 4 gnd
rlabel metal3 s 9182 4385 9280 4483 4 vdd
rlabel metal3 s 6698 5545 6796 5643 4 gnd
rlabel metal3 s 9194 5545 9292 5643 4 gnd
rlabel metal3 s 2954 5545 3052 5643 4 gnd
rlabel metal3 s 14174 4385 14272 4483 4 vdd
rlabel metal3 s 3024 3611 3122 3709 4 gnd
rlabel metal3 s 16682 5545 16780 5643 4 gnd
rlabel metal3 s 5450 5545 5548 5643 4 gnd
rlabel metal3 s 8016 3611 8114 3709 4 gnd
rlabel metal3 s 20426 5545 20524 5643 4 gnd
rlabel metal3 s 3197 1862 3295 1960 4 gnd
rlabel metal3 s 15434 5545 15532 5643 4 gnd
rlabel metal3 s 10512 3611 10610 3709 4 gnd
rlabel metal3 s 15677 1862 15775 1960 4 gnd
rlabel metal3 s 13008 3611 13106 3709 4 gnd
rlabel metal3 s 11760 3611 11858 3709 4 gnd
rlabel metal3 s 17930 5545 18028 5643 4 gnd
rlabel metal3 s 12750 313 12848 411 4 vdd
rlabel metal3 s 4014 313 4112 411 4 vdd
rlabel metal3 s 3628 313 3726 411 4 vdd
rlabel metal3 s 15246 313 15344 411 4 vdd
rlabel metal3 s 20238 313 20336 411 4 vdd
rlabel metal3 s 10254 313 10352 411 4 vdd
rlabel metal3 s 14860 313 14958 411 4 vdd
rlabel metal3 s 13998 313 14096 411 4 vdd
rlabel metal3 s 17356 313 17454 411 4 vdd
rlabel metal3 s 13612 313 13710 411 4 vdd
rlabel metal3 s 2766 313 2864 411 4 vdd
rlabel metal3 s 12364 313 12462 411 4 vdd
rlabel metal3 s 21486 313 21584 411 4 vdd
rlabel metal3 s 16108 313 16206 411 4 vdd
rlabel metal3 s 6124 313 6222 411 4 vdd
rlabel metal3 s 18604 313 18702 411 4 vdd
rlabel metal3 s 7758 313 7856 411 4 vdd
rlabel metal3 s 16494 313 16592 411 4 vdd
rlabel metal3 s 8620 313 8718 411 4 vdd
rlabel metal3 s 21100 313 21198 411 4 vdd
rlabel metal3 s 6510 313 6608 411 4 vdd
rlabel metal3 s 4876 313 4974 411 4 vdd
rlabel metal3 s 17742 313 17840 411 4 vdd
rlabel metal3 s 2380 313 2478 411 4 vdd
rlabel metal3 s 7372 313 7470 411 4 vdd
rlabel metal3 s 9868 313 9966 411 4 vdd
rlabel metal3 s 18990 313 19088 411 4 vdd
rlabel metal3 s 9006 313 9104 411 4 vdd
rlabel metal3 s 5262 313 5360 411 4 vdd
rlabel metal3 s 19852 313 19950 411 4 vdd
rlabel metal3 s 11116 313 11214 411 4 vdd
rlabel metal3 s 1518 313 1616 411 4 vdd
rlabel metal3 s 11502 313 11600 411 4 vdd
rlabel metal3 s 32718 313 32816 411 4 vdd
rlabel metal3 s 27726 313 27824 411 4 vdd
rlabel metal3 s 30222 313 30320 411 4 vdd
rlabel metal3 s 37324 313 37422 411 4 vdd
rlabel metal3 s 39820 313 39918 411 4 vdd
rlabel metal3 s 24844 313 24942 411 4 vdd
rlabel metal3 s 38572 313 38670 411 4 vdd
rlabel metal3 s 36076 313 36174 411 4 vdd
rlabel metal3 s 40206 313 40304 411 4 vdd
rlabel metal3 s 29836 313 29934 411 4 vdd
rlabel metal3 s 28588 313 28686 411 4 vdd
rlabel metal3 s 33966 313 34064 411 4 vdd
rlabel metal3 s 22348 313 22446 411 4 vdd
rlabel metal3 s 35214 313 35312 411 4 vdd
rlabel metal3 s 37710 313 37808 411 4 vdd
rlabel metal3 s 41454 313 41552 411 4 vdd
rlabel metal3 s 23982 313 24080 411 4 vdd
rlabel metal3 s 26478 313 26576 411 4 vdd
rlabel metal3 s 32332 313 32430 411 4 vdd
rlabel metal3 s 36462 313 36560 411 4 vdd
rlabel metal3 s 28974 313 29072 411 4 vdd
rlabel metal3 s 38958 313 39056 411 4 vdd
rlabel metal3 s 31470 313 31568 411 4 vdd
rlabel metal3 s 41068 313 41166 411 4 vdd
rlabel metal3 s 31084 313 31182 411 4 vdd
rlabel metal3 s 33580 313 33678 411 4 vdd
rlabel metal3 s 34828 313 34926 411 4 vdd
rlabel metal3 s 25230 313 25328 411 4 vdd
rlabel metal3 s 22734 313 22832 411 4 vdd
rlabel metal3 s 27340 313 27438 411 4 vdd
rlabel metal3 s 26092 313 26190 411 4 vdd
rlabel metal3 s 23596 313 23694 411 4 vdd
rlabel metal1 s 22694 5448 22740 5702 4 dout_17
rlabel metal1 s 23942 5448 23988 5702 4 dout_18
rlabel metal1 s 25190 5448 25236 5702 4 dout_19
rlabel metal1 s 26438 5448 26484 5702 4 dout_20
rlabel metal1 s 27686 5448 27732 5702 4 dout_21
rlabel metal1 s 28934 5448 28980 5702 4 dout_22
rlabel metal1 s 30182 5448 30228 5702 4 dout_23
rlabel metal1 s 31430 5448 31476 5702 4 dout_24
rlabel metal1 s 32678 5448 32724 5702 4 dout_25
rlabel metal1 s 33926 5448 33972 5702 4 dout_26
rlabel metal1 s 35174 5448 35220 5702 4 dout_27
rlabel metal1 s 36422 5448 36468 5702 4 dout_28
rlabel metal1 s 37670 5448 37716 5702 4 dout_29
rlabel metal1 s 38918 5448 38964 5702 4 dout_30
rlabel metal1 s 40166 5448 40212 5702 4 dout_31
rlabel metal1 s 20198 5448 20244 5702 4 dout_15
rlabel metal1 s 21446 5448 21492 5702 4 dout_16
rlabel metal1 s 1478 5448 1524 5702 4 dout_0
rlabel metal1 s 2726 5448 2772 5702 4 dout_1
rlabel metal1 s 3974 5448 4020 5702 4 dout_2
rlabel metal1 s 5222 5448 5268 5702 4 dout_3
rlabel metal1 s 6470 5448 6516 5702 4 dout_4
rlabel metal1 s 7718 5448 7764 5702 4 dout_5
rlabel metal1 s 8966 5448 9012 5702 4 dout_6
rlabel metal1 s 10214 5448 10260 5702 4 dout_7
rlabel metal1 s 11462 5448 11508 5702 4 dout_8
rlabel metal1 s 12710 5448 12756 5702 4 dout_9
rlabel metal1 s 13958 5448 14004 5702 4 dout_10
rlabel metal1 s 15206 5448 15252 5702 4 dout_11
rlabel metal1 s 16454 5448 16500 5702 4 dout_12
rlabel metal1 s 17702 5448 17748 5702 4 dout_13
rlabel metal1 s 18950 5448 18996 5702 4 dout_14
rlabel metal1 s 1440 252 1468 1006 4 bl_0
rlabel metal1 s 1904 252 1932 1006 4 br_0
rlabel metal1 s 2528 252 2556 1006 4 bl_1
rlabel metal1 s 2064 252 2092 1006 4 br_1
rlabel metal1 s 2688 252 2716 1006 4 bl_2
rlabel metal1 s 3152 252 3180 1006 4 br_2
rlabel metal1 s 3776 252 3804 1006 4 bl_3
rlabel metal1 s 3312 252 3340 1006 4 br_3
rlabel metal1 s 3936 252 3964 1006 4 bl_4
rlabel metal1 s 4400 252 4428 1006 4 br_4
rlabel metal1 s 5024 252 5052 1006 4 bl_5
rlabel metal1 s 4560 252 4588 1006 4 br_5
rlabel metal1 s 5184 252 5212 1006 4 bl_6
rlabel metal1 s 5648 252 5676 1006 4 br_6
rlabel metal1 s 6272 252 6300 1006 4 bl_7
rlabel metal1 s 5808 252 5836 1006 4 br_7
rlabel metal1 s 6432 252 6460 1006 4 bl_8
rlabel metal1 s 6896 252 6924 1006 4 br_8
rlabel metal1 s 7520 252 7548 1006 4 bl_9
rlabel metal1 s 7056 252 7084 1006 4 br_9
rlabel metal1 s 7680 252 7708 1006 4 bl_10
rlabel metal1 s 8144 252 8172 1006 4 br_10
rlabel metal1 s 8768 252 8796 1006 4 bl_11
rlabel metal1 s 8304 252 8332 1006 4 br_11
rlabel metal1 s 8928 252 8956 1006 4 bl_12
rlabel metal1 s 9392 252 9420 1006 4 br_12
rlabel metal1 s 10016 252 10044 1006 4 bl_13
rlabel metal1 s 9552 252 9580 1006 4 br_13
rlabel metal1 s 10176 252 10204 1006 4 bl_14
rlabel metal1 s 10640 252 10668 1006 4 br_14
rlabel metal1 s 11264 252 11292 1006 4 bl_15
rlabel metal1 s 10800 252 10828 1006 4 br_15
rlabel metal1 s 11424 252 11452 1006 4 bl_16
rlabel metal1 s 11888 252 11916 1006 4 br_16
rlabel metal1 s 12512 252 12540 1006 4 bl_17
rlabel metal1 s 12048 252 12076 1006 4 br_17
rlabel metal1 s 12672 252 12700 1006 4 bl_18
rlabel metal1 s 13136 252 13164 1006 4 br_18
rlabel metal1 s 13760 252 13788 1006 4 bl_19
rlabel metal1 s 13296 252 13324 1006 4 br_19
rlabel metal1 s 13920 252 13948 1006 4 bl_20
rlabel metal1 s 14384 252 14412 1006 4 br_20
rlabel metal1 s 15008 252 15036 1006 4 bl_21
rlabel metal1 s 14544 252 14572 1006 4 br_21
rlabel metal1 s 15168 252 15196 1006 4 bl_22
rlabel metal1 s 15632 252 15660 1006 4 br_22
rlabel metal1 s 16256 252 16284 1006 4 bl_23
rlabel metal1 s 15792 252 15820 1006 4 br_23
rlabel metal1 s 16416 252 16444 1006 4 bl_24
rlabel metal1 s 16880 252 16908 1006 4 br_24
rlabel metal1 s 17504 252 17532 1006 4 bl_25
rlabel metal1 s 17040 252 17068 1006 4 br_25
rlabel metal1 s 17664 252 17692 1006 4 bl_26
rlabel metal1 s 18128 252 18156 1006 4 br_26
rlabel metal1 s 18752 252 18780 1006 4 bl_27
rlabel metal1 s 18288 252 18316 1006 4 br_27
rlabel metal1 s 18912 252 18940 1006 4 bl_28
rlabel metal1 s 19376 252 19404 1006 4 br_28
rlabel metal1 s 20000 252 20028 1006 4 bl_29
rlabel metal1 s 19536 252 19564 1006 4 br_29
rlabel metal1 s 20160 252 20188 1006 4 bl_30
rlabel metal1 s 20624 252 20652 1006 4 br_30
rlabel metal1 s 21248 252 21276 1006 4 bl_31
rlabel metal1 s 20784 252 20812 1006 4 br_31
rlabel metal1 s 21408 252 21436 1006 4 bl_32
rlabel metal1 s 41840 252 41868 1006 4 rbl_br
rlabel metal1 s 41376 252 41404 1006 4 rbl_bl
rlabel metal1 s 21872 252 21900 1006 4 br_32
rlabel metal1 s 22496 252 22524 1006 4 bl_33
rlabel metal1 s 22032 252 22060 1006 4 br_33
rlabel metal1 s 22656 252 22684 1006 4 bl_34
rlabel metal1 s 23120 252 23148 1006 4 br_34
rlabel metal1 s 23744 252 23772 1006 4 bl_35
rlabel metal1 s 23280 252 23308 1006 4 br_35
rlabel metal1 s 23904 252 23932 1006 4 bl_36
rlabel metal1 s 24368 252 24396 1006 4 br_36
rlabel metal1 s 24992 252 25020 1006 4 bl_37
rlabel metal1 s 24528 252 24556 1006 4 br_37
rlabel metal1 s 25152 252 25180 1006 4 bl_38
rlabel metal1 s 25616 252 25644 1006 4 br_38
rlabel metal1 s 26240 252 26268 1006 4 bl_39
rlabel metal1 s 25776 252 25804 1006 4 br_39
rlabel metal1 s 26400 252 26428 1006 4 bl_40
rlabel metal1 s 26864 252 26892 1006 4 br_40
rlabel metal1 s 27488 252 27516 1006 4 bl_41
rlabel metal1 s 27024 252 27052 1006 4 br_41
rlabel metal1 s 27648 252 27676 1006 4 bl_42
rlabel metal1 s 28112 252 28140 1006 4 br_42
rlabel metal1 s 28736 252 28764 1006 4 bl_43
rlabel metal1 s 28272 252 28300 1006 4 br_43
rlabel metal1 s 28896 252 28924 1006 4 bl_44
rlabel metal1 s 29360 252 29388 1006 4 br_44
rlabel metal1 s 29984 252 30012 1006 4 bl_45
rlabel metal1 s 29520 252 29548 1006 4 br_45
rlabel metal1 s 30144 252 30172 1006 4 bl_46
rlabel metal1 s 30608 252 30636 1006 4 br_46
rlabel metal1 s 31232 252 31260 1006 4 bl_47
rlabel metal1 s 30768 252 30796 1006 4 br_47
rlabel metal1 s 31392 252 31420 1006 4 bl_48
rlabel metal1 s 31856 252 31884 1006 4 br_48
rlabel metal1 s 32480 252 32508 1006 4 bl_49
rlabel metal1 s 32016 252 32044 1006 4 br_49
rlabel metal1 s 32640 252 32668 1006 4 bl_50
rlabel metal1 s 33104 252 33132 1006 4 br_50
rlabel metal1 s 33728 252 33756 1006 4 bl_51
rlabel metal1 s 33264 252 33292 1006 4 br_51
rlabel metal1 s 33888 252 33916 1006 4 bl_52
rlabel metal1 s 34352 252 34380 1006 4 br_52
rlabel metal1 s 34976 252 35004 1006 4 bl_53
rlabel metal1 s 34512 252 34540 1006 4 br_53
rlabel metal1 s 35136 252 35164 1006 4 bl_54
rlabel metal1 s 35600 252 35628 1006 4 br_54
rlabel metal1 s 36224 252 36252 1006 4 bl_55
rlabel metal1 s 35760 252 35788 1006 4 br_55
rlabel metal1 s 36384 252 36412 1006 4 bl_56
rlabel metal1 s 36848 252 36876 1006 4 br_56
rlabel metal1 s 37472 252 37500 1006 4 bl_57
rlabel metal1 s 37008 252 37036 1006 4 br_57
rlabel metal1 s 37632 252 37660 1006 4 bl_58
rlabel metal1 s 38096 252 38124 1006 4 br_58
rlabel metal1 s 38720 252 38748 1006 4 bl_59
rlabel metal1 s 38256 252 38284 1006 4 br_59
rlabel metal1 s 38880 252 38908 1006 4 bl_60
rlabel metal1 s 39344 252 39372 1006 4 br_60
rlabel metal1 s 39968 252 39996 1006 4 bl_61
rlabel metal1 s 39504 252 39532 1006 4 br_61
rlabel metal1 s 40128 252 40156 1006 4 bl_62
rlabel metal1 s 40592 252 40620 1006 4 br_62
rlabel metal1 s 41216 252 41244 1006 4 bl_63
rlabel metal1 s 40752 252 40780 1006 4 br_63
<< properties >>
string FIXED_BBOX 0 0 41934 5702
string GDS_END 6801034
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 6670848
<< end >>
