magic
tech sky130B
magscale 1 2
timestamp 1676037725
use sky130_fd_pr__via_l1m1__example_55959141808683  sky130_fd_pr__via_l1m1__example_55959141808683_0
timestamp 1676037725
transform 1 0 61 0 1 139
box 0 0 1 1
<< properties >>
string GDS_END 8041566
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8028468
<< end >>
