/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.ref/sky130_fd_io/lef/sky130_fd_io.lef