/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/xschem/xschem_verilog_import/audiodac.spice