magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
rect 78 0 114 395
rect 150 0 186 395
rect 294 0 330 395
rect 366 0 402 395
rect 846 0 882 395
rect 918 0 954 395
rect 1062 0 1098 395
rect 1134 0 1170 395
rect 1326 0 1362 395
rect 1398 0 1434 395
rect 1542 0 1578 395
rect 1614 0 1650 395
rect 2094 0 2130 395
rect 2166 0 2202 395
rect 2310 0 2346 395
rect 2382 0 2418 395
rect 2574 0 2610 395
rect 2646 0 2682 395
rect 2790 0 2826 395
rect 2862 0 2898 395
rect 3342 0 3378 395
rect 3414 0 3450 395
rect 3558 0 3594 395
rect 3630 0 3666 395
rect 3822 0 3858 395
rect 3894 0 3930 395
rect 4038 0 4074 395
rect 4110 0 4146 395
rect 4590 0 4626 395
rect 4662 0 4698 395
rect 4806 0 4842 395
rect 4878 0 4914 395
rect 5070 0 5106 395
rect 5142 0 5178 395
rect 5286 0 5322 395
rect 5358 0 5394 395
rect 5838 0 5874 395
rect 5910 0 5946 395
rect 6054 0 6090 395
rect 6126 0 6162 395
rect 6318 0 6354 395
rect 6390 0 6426 395
rect 6534 0 6570 395
rect 6606 0 6642 395
rect 7086 0 7122 395
rect 7158 0 7194 395
rect 7302 0 7338 395
rect 7374 0 7410 395
rect 7566 0 7602 395
rect 7638 0 7674 395
rect 7782 0 7818 395
rect 7854 0 7890 395
rect 8334 0 8370 395
rect 8406 0 8442 395
rect 8550 0 8586 395
rect 8622 0 8658 395
rect 8814 0 8850 395
rect 8886 0 8922 395
rect 9030 0 9066 395
rect 9102 0 9138 395
rect 9582 0 9618 395
rect 9654 0 9690 395
rect 9798 0 9834 395
rect 9870 0 9906 395
rect 10062 0 10098 395
rect 10134 0 10170 395
rect 10278 0 10314 395
rect 10350 0 10386 395
rect 10830 0 10866 395
rect 10902 0 10938 395
rect 11046 0 11082 395
rect 11118 0 11154 395
rect 11310 0 11346 395
rect 11382 0 11418 395
rect 11526 0 11562 395
rect 11598 0 11634 395
rect 12078 0 12114 395
rect 12150 0 12186 395
rect 12294 0 12330 395
rect 12366 0 12402 395
rect 12558 0 12594 395
rect 12630 0 12666 395
rect 12774 0 12810 395
rect 12846 0 12882 395
rect 13326 0 13362 395
rect 13398 0 13434 395
rect 13542 0 13578 395
rect 13614 0 13650 395
rect 13806 0 13842 395
rect 13878 0 13914 395
rect 14022 0 14058 395
rect 14094 0 14130 395
rect 14574 0 14610 395
rect 14646 0 14682 395
rect 14790 0 14826 395
rect 14862 0 14898 395
rect 15054 0 15090 395
rect 15126 0 15162 395
rect 15270 0 15306 395
rect 15342 0 15378 395
rect 15822 0 15858 395
rect 15894 0 15930 395
rect 16038 0 16074 395
rect 16110 0 16146 395
rect 16302 0 16338 395
rect 16374 0 16410 395
rect 16518 0 16554 395
rect 16590 0 16626 395
rect 17070 0 17106 395
rect 17142 0 17178 395
rect 17286 0 17322 395
rect 17358 0 17394 395
rect 17550 0 17586 395
rect 17622 0 17658 395
rect 17766 0 17802 395
rect 17838 0 17874 395
rect 18318 0 18354 395
rect 18390 0 18426 395
rect 18534 0 18570 395
rect 18606 0 18642 395
rect 18798 0 18834 395
rect 18870 0 18906 395
rect 19014 0 19050 395
rect 19086 0 19122 395
rect 19566 0 19602 395
rect 19638 0 19674 395
rect 19782 0 19818 395
rect 19854 0 19890 395
rect 20046 0 20082 395
rect 20118 0 20154 395
rect 20262 0 20298 395
rect 20334 0 20370 395
rect 20814 0 20850 395
rect 20886 0 20922 395
rect 21030 0 21066 395
rect 21102 0 21138 395
rect 21294 0 21330 395
rect 21366 0 21402 395
rect 21510 0 21546 395
rect 21582 0 21618 395
rect 22062 0 22098 395
rect 22134 0 22170 395
rect 22278 0 22314 395
rect 22350 0 22386 395
rect 22542 0 22578 395
rect 22614 0 22650 395
rect 22758 0 22794 395
rect 22830 0 22866 395
rect 23310 0 23346 395
rect 23382 0 23418 395
rect 23526 0 23562 395
rect 23598 0 23634 395
rect 23790 0 23826 395
rect 23862 0 23898 395
rect 24006 0 24042 395
rect 24078 0 24114 395
rect 24558 0 24594 395
rect 24630 0 24666 395
rect 24774 0 24810 395
rect 24846 0 24882 395
rect 25038 0 25074 395
rect 25110 0 25146 395
rect 25254 0 25290 395
rect 25326 0 25362 395
rect 25806 0 25842 395
rect 25878 0 25914 395
rect 26022 0 26058 395
rect 26094 0 26130 395
rect 26286 0 26322 395
rect 26358 0 26394 395
rect 26502 0 26538 395
rect 26574 0 26610 395
rect 27054 0 27090 395
rect 27126 0 27162 395
rect 27270 0 27306 395
rect 27342 0 27378 395
rect 27534 0 27570 395
rect 27606 0 27642 395
rect 27750 0 27786 395
rect 27822 0 27858 395
rect 28302 0 28338 395
rect 28374 0 28410 395
rect 28518 0 28554 395
rect 28590 0 28626 395
rect 28782 0 28818 395
rect 28854 0 28890 395
rect 28998 0 29034 395
rect 29070 0 29106 395
rect 29550 0 29586 395
rect 29622 0 29658 395
rect 29766 0 29802 395
rect 29838 0 29874 395
rect 30030 0 30066 395
rect 30102 0 30138 395
rect 30246 0 30282 395
rect 30318 0 30354 395
rect 30798 0 30834 395
rect 30870 0 30906 395
rect 31014 0 31050 395
rect 31086 0 31122 395
rect 31278 0 31314 395
rect 31350 0 31386 395
rect 31494 0 31530 395
rect 31566 0 31602 395
rect 32046 0 32082 395
rect 32118 0 32154 395
rect 32262 0 32298 395
rect 32334 0 32370 395
rect 32526 0 32562 395
rect 32598 0 32634 395
rect 32742 0 32778 395
rect 32814 0 32850 395
rect 33294 0 33330 395
rect 33366 0 33402 395
rect 33510 0 33546 395
rect 33582 0 33618 395
rect 33774 0 33810 395
rect 33846 0 33882 395
rect 33990 0 34026 395
rect 34062 0 34098 395
rect 34542 0 34578 395
rect 34614 0 34650 395
rect 34758 0 34794 395
rect 34830 0 34866 395
rect 35022 0 35058 395
rect 35094 0 35130 395
rect 35238 0 35274 395
rect 35310 0 35346 395
rect 35790 0 35826 395
rect 35862 0 35898 395
rect 36006 0 36042 395
rect 36078 0 36114 395
rect 36270 0 36306 395
rect 36342 0 36378 395
rect 36486 0 36522 395
rect 36558 0 36594 395
rect 37038 0 37074 395
rect 37110 0 37146 395
rect 37254 0 37290 395
rect 37326 0 37362 395
rect 37518 0 37554 395
rect 37590 0 37626 395
rect 37734 0 37770 395
rect 37806 0 37842 395
rect 38286 0 38322 395
rect 38358 0 38394 395
rect 38502 0 38538 395
rect 38574 0 38610 395
rect 38766 0 38802 395
rect 38838 0 38874 395
rect 38982 0 39018 395
rect 39054 0 39090 395
rect 39534 0 39570 395
rect 39606 0 39642 395
rect 39750 0 39786 395
rect 39822 0 39858 395
rect 40014 0 40050 395
rect 40086 0 40122 395
rect 40230 0 40266 395
rect 40302 0 40338 395
rect 40782 0 40818 395
rect 40854 0 40890 395
rect 40998 0 41034 395
rect 41070 0 41106 395
rect 41262 0 41298 395
rect 41334 0 41370 395
rect 41478 0 41514 395
rect 41550 0 41586 395
rect 42030 0 42066 395
rect 42102 0 42138 395
rect 42246 0 42282 395
rect 42318 0 42354 395
rect 42510 0 42546 395
rect 42582 0 42618 395
rect 42726 0 42762 395
rect 42798 0 42834 395
rect 43278 0 43314 395
rect 43350 0 43386 395
rect 43494 0 43530 395
rect 43566 0 43602 395
rect 43758 0 43794 395
rect 43830 0 43866 395
rect 43974 0 44010 395
rect 44046 0 44082 395
rect 44526 0 44562 395
rect 44598 0 44634 395
rect 44742 0 44778 395
rect 44814 0 44850 395
rect 45006 0 45042 395
rect 45078 0 45114 395
rect 45222 0 45258 395
rect 45294 0 45330 395
rect 45774 0 45810 395
rect 45846 0 45882 395
rect 45990 0 46026 395
rect 46062 0 46098 395
rect 46254 0 46290 395
rect 46326 0 46362 395
rect 46470 0 46506 395
rect 46542 0 46578 395
rect 47022 0 47058 395
rect 47094 0 47130 395
rect 47238 0 47274 395
rect 47310 0 47346 395
rect 47502 0 47538 395
rect 47574 0 47610 395
rect 47718 0 47754 395
rect 47790 0 47826 395
rect 48270 0 48306 395
rect 48342 0 48378 395
rect 48486 0 48522 395
rect 48558 0 48594 395
rect 48750 0 48786 395
rect 48822 0 48858 395
rect 48966 0 49002 395
rect 49038 0 49074 395
rect 49518 0 49554 395
rect 49590 0 49626 395
rect 49734 0 49770 395
rect 49806 0 49842 395
rect 49998 0 50034 395
rect 50070 0 50106 395
rect 50214 0 50250 395
rect 50286 0 50322 395
rect 50766 0 50802 395
rect 50838 0 50874 395
rect 50982 0 51018 395
rect 51054 0 51090 395
rect 51246 0 51282 395
rect 51318 0 51354 395
rect 51462 0 51498 395
rect 51534 0 51570 395
rect 52014 0 52050 395
rect 52086 0 52122 395
rect 52230 0 52266 395
rect 52302 0 52338 395
rect 52494 0 52530 395
rect 52566 0 52602 395
rect 52710 0 52746 395
rect 52782 0 52818 395
rect 53262 0 53298 395
rect 53334 0 53370 395
rect 53478 0 53514 395
rect 53550 0 53586 395
rect 53742 0 53778 395
rect 53814 0 53850 395
rect 53958 0 53994 395
rect 54030 0 54066 395
rect 54510 0 54546 395
rect 54582 0 54618 395
rect 54726 0 54762 395
rect 54798 0 54834 395
rect 54990 0 55026 395
rect 55062 0 55098 395
rect 55206 0 55242 395
rect 55278 0 55314 395
rect 55758 0 55794 395
rect 55830 0 55866 395
rect 55974 0 56010 395
rect 56046 0 56082 395
rect 56238 0 56274 395
rect 56310 0 56346 395
rect 56454 0 56490 395
rect 56526 0 56562 395
rect 57006 0 57042 395
rect 57078 0 57114 395
rect 57222 0 57258 395
rect 57294 0 57330 395
rect 57486 0 57522 395
rect 57558 0 57594 395
rect 57702 0 57738 395
rect 57774 0 57810 395
rect 58254 0 58290 395
rect 58326 0 58362 395
rect 58470 0 58506 395
rect 58542 0 58578 395
rect 58734 0 58770 395
rect 58806 0 58842 395
rect 58950 0 58986 395
rect 59022 0 59058 395
rect 59502 0 59538 395
rect 59574 0 59610 395
rect 59718 0 59754 395
rect 59790 0 59826 395
rect 59982 0 60018 395
rect 60054 0 60090 395
rect 60198 0 60234 395
rect 60270 0 60306 395
rect 60750 0 60786 395
rect 60822 0 60858 395
rect 60966 0 61002 395
rect 61038 0 61074 395
rect 61230 0 61266 395
rect 61302 0 61338 395
rect 61446 0 61482 395
rect 61518 0 61554 395
rect 61998 0 62034 395
rect 62070 0 62106 395
rect 62214 0 62250 395
rect 62286 0 62322 395
rect 62478 0 62514 395
rect 62550 0 62586 395
rect 62694 0 62730 395
rect 62766 0 62802 395
rect 63246 0 63282 395
rect 63318 0 63354 395
rect 63462 0 63498 395
rect 63534 0 63570 395
rect 63726 0 63762 395
rect 63798 0 63834 395
rect 63942 0 63978 395
rect 64014 0 64050 395
rect 64494 0 64530 395
rect 64566 0 64602 395
rect 64710 0 64746 395
rect 64782 0 64818 395
rect 64974 0 65010 395
rect 65046 0 65082 395
rect 65190 0 65226 395
rect 65262 0 65298 395
rect 65742 0 65778 395
rect 65814 0 65850 395
rect 65958 0 65994 395
rect 66030 0 66066 395
rect 66222 0 66258 395
rect 66294 0 66330 395
rect 66438 0 66474 395
rect 66510 0 66546 395
rect 66990 0 67026 395
rect 67062 0 67098 395
rect 67206 0 67242 395
rect 67278 0 67314 395
rect 67470 0 67506 395
rect 67542 0 67578 395
rect 67686 0 67722 395
rect 67758 0 67794 395
rect 68238 0 68274 395
rect 68310 0 68346 395
rect 68454 0 68490 395
rect 68526 0 68562 395
rect 68718 0 68754 395
rect 68790 0 68826 395
rect 68934 0 68970 395
rect 69006 0 69042 395
rect 69486 0 69522 395
rect 69558 0 69594 395
rect 69702 0 69738 395
rect 69774 0 69810 395
rect 69966 0 70002 395
rect 70038 0 70074 395
rect 70182 0 70218 395
rect 70254 0 70290 395
rect 70734 0 70770 395
rect 70806 0 70842 395
rect 70950 0 70986 395
rect 71022 0 71058 395
rect 71214 0 71250 395
rect 71286 0 71322 395
rect 71430 0 71466 395
rect 71502 0 71538 395
rect 71982 0 72018 395
rect 72054 0 72090 395
rect 72198 0 72234 395
rect 72270 0 72306 395
rect 72462 0 72498 395
rect 72534 0 72570 395
rect 72678 0 72714 395
rect 72750 0 72786 395
rect 73230 0 73266 395
rect 73302 0 73338 395
rect 73446 0 73482 395
rect 73518 0 73554 395
rect 73710 0 73746 395
rect 73782 0 73818 395
rect 73926 0 73962 395
rect 73998 0 74034 395
rect 74478 0 74514 395
rect 74550 0 74586 395
rect 74694 0 74730 395
rect 74766 0 74802 395
rect 74958 0 74994 395
rect 75030 0 75066 395
rect 75174 0 75210 395
rect 75246 0 75282 395
rect 75726 0 75762 395
rect 75798 0 75834 395
rect 75942 0 75978 395
rect 76014 0 76050 395
rect 76206 0 76242 395
rect 76278 0 76314 395
rect 76422 0 76458 395
rect 76494 0 76530 395
rect 76974 0 77010 395
rect 77046 0 77082 395
rect 77190 0 77226 395
rect 77262 0 77298 395
rect 77454 0 77490 395
rect 77526 0 77562 395
rect 77670 0 77706 395
rect 77742 0 77778 395
rect 78222 0 78258 395
rect 78294 0 78330 395
rect 78438 0 78474 395
rect 78510 0 78546 395
rect 78702 0 78738 395
rect 78774 0 78810 395
rect 78918 0 78954 395
rect 78990 0 79026 395
rect 79470 0 79506 395
rect 79542 0 79578 395
rect 79686 0 79722 395
rect 79758 0 79794 395
<< metal2 >>
rect 284 257 340 266
rect 284 192 340 201
rect 908 257 964 266
rect 908 192 964 201
rect 1532 257 1588 266
rect 1532 192 1588 201
rect 2156 257 2212 266
rect 2156 192 2212 201
rect 2780 257 2836 266
rect 2780 192 2836 201
rect 3404 257 3460 266
rect 3404 192 3460 201
rect 4028 257 4084 266
rect 4028 192 4084 201
rect 4652 257 4708 266
rect 4652 192 4708 201
rect 5276 257 5332 266
rect 5276 192 5332 201
rect 5900 257 5956 266
rect 5900 192 5956 201
rect 6524 257 6580 266
rect 6524 192 6580 201
rect 7148 257 7204 266
rect 7148 192 7204 201
rect 7772 257 7828 266
rect 7772 192 7828 201
rect 8396 257 8452 266
rect 8396 192 8452 201
rect 9020 257 9076 266
rect 9020 192 9076 201
rect 9644 257 9700 266
rect 9644 192 9700 201
rect 10268 257 10324 266
rect 10268 192 10324 201
rect 10892 257 10948 266
rect 10892 192 10948 201
rect 11516 257 11572 266
rect 11516 192 11572 201
rect 12140 257 12196 266
rect 12140 192 12196 201
rect 12764 257 12820 266
rect 12764 192 12820 201
rect 13388 257 13444 266
rect 13388 192 13444 201
rect 14012 257 14068 266
rect 14012 192 14068 201
rect 14636 257 14692 266
rect 14636 192 14692 201
rect 15260 257 15316 266
rect 15260 192 15316 201
rect 15884 257 15940 266
rect 15884 192 15940 201
rect 16508 257 16564 266
rect 16508 192 16564 201
rect 17132 257 17188 266
rect 17132 192 17188 201
rect 17756 257 17812 266
rect 17756 192 17812 201
rect 18380 257 18436 266
rect 18380 192 18436 201
rect 19004 257 19060 266
rect 19004 192 19060 201
rect 19628 257 19684 266
rect 19628 192 19684 201
rect 20252 257 20308 266
rect 20252 192 20308 201
rect 20876 257 20932 266
rect 20876 192 20932 201
rect 21500 257 21556 266
rect 21500 192 21556 201
rect 22124 257 22180 266
rect 22124 192 22180 201
rect 22748 257 22804 266
rect 22748 192 22804 201
rect 23372 257 23428 266
rect 23372 192 23428 201
rect 23996 257 24052 266
rect 23996 192 24052 201
rect 24620 257 24676 266
rect 24620 192 24676 201
rect 25244 257 25300 266
rect 25244 192 25300 201
rect 25868 257 25924 266
rect 25868 192 25924 201
rect 26492 257 26548 266
rect 26492 192 26548 201
rect 27116 257 27172 266
rect 27116 192 27172 201
rect 27740 257 27796 266
rect 27740 192 27796 201
rect 28364 257 28420 266
rect 28364 192 28420 201
rect 28988 257 29044 266
rect 28988 192 29044 201
rect 29612 257 29668 266
rect 29612 192 29668 201
rect 30236 257 30292 266
rect 30236 192 30292 201
rect 30860 257 30916 266
rect 30860 192 30916 201
rect 31484 257 31540 266
rect 31484 192 31540 201
rect 32108 257 32164 266
rect 32108 192 32164 201
rect 32732 257 32788 266
rect 32732 192 32788 201
rect 33356 257 33412 266
rect 33356 192 33412 201
rect 33980 257 34036 266
rect 33980 192 34036 201
rect 34604 257 34660 266
rect 34604 192 34660 201
rect 35228 257 35284 266
rect 35228 192 35284 201
rect 35852 257 35908 266
rect 35852 192 35908 201
rect 36476 257 36532 266
rect 36476 192 36532 201
rect 37100 257 37156 266
rect 37100 192 37156 201
rect 37724 257 37780 266
rect 37724 192 37780 201
rect 38348 257 38404 266
rect 38348 192 38404 201
rect 38972 257 39028 266
rect 38972 192 39028 201
rect 39596 257 39652 266
rect 39596 192 39652 201
rect 40220 257 40276 266
rect 40220 192 40276 201
rect 40844 257 40900 266
rect 40844 192 40900 201
rect 41468 257 41524 266
rect 41468 192 41524 201
rect 42092 257 42148 266
rect 42092 192 42148 201
rect 42716 257 42772 266
rect 42716 192 42772 201
rect 43340 257 43396 266
rect 43340 192 43396 201
rect 43964 257 44020 266
rect 43964 192 44020 201
rect 44588 257 44644 266
rect 44588 192 44644 201
rect 45212 257 45268 266
rect 45212 192 45268 201
rect 45836 257 45892 266
rect 45836 192 45892 201
rect 46460 257 46516 266
rect 46460 192 46516 201
rect 47084 257 47140 266
rect 47084 192 47140 201
rect 47708 257 47764 266
rect 47708 192 47764 201
rect 48332 257 48388 266
rect 48332 192 48388 201
rect 48956 257 49012 266
rect 48956 192 49012 201
rect 49580 257 49636 266
rect 49580 192 49636 201
rect 50204 257 50260 266
rect 50204 192 50260 201
rect 50828 257 50884 266
rect 50828 192 50884 201
rect 51452 257 51508 266
rect 51452 192 51508 201
rect 52076 257 52132 266
rect 52076 192 52132 201
rect 52700 257 52756 266
rect 52700 192 52756 201
rect 53324 257 53380 266
rect 53324 192 53380 201
rect 53948 257 54004 266
rect 53948 192 54004 201
rect 54572 257 54628 266
rect 54572 192 54628 201
rect 55196 257 55252 266
rect 55196 192 55252 201
rect 55820 257 55876 266
rect 55820 192 55876 201
rect 56444 257 56500 266
rect 56444 192 56500 201
rect 57068 257 57124 266
rect 57068 192 57124 201
rect 57692 257 57748 266
rect 57692 192 57748 201
rect 58316 257 58372 266
rect 58316 192 58372 201
rect 58940 257 58996 266
rect 58940 192 58996 201
rect 59564 257 59620 266
rect 59564 192 59620 201
rect 60188 257 60244 266
rect 60188 192 60244 201
rect 60812 257 60868 266
rect 60812 192 60868 201
rect 61436 257 61492 266
rect 61436 192 61492 201
rect 62060 257 62116 266
rect 62060 192 62116 201
rect 62684 257 62740 266
rect 62684 192 62740 201
rect 63308 257 63364 266
rect 63308 192 63364 201
rect 63932 257 63988 266
rect 63932 192 63988 201
rect 64556 257 64612 266
rect 64556 192 64612 201
rect 65180 257 65236 266
rect 65180 192 65236 201
rect 65804 257 65860 266
rect 65804 192 65860 201
rect 66428 257 66484 266
rect 66428 192 66484 201
rect 67052 257 67108 266
rect 67052 192 67108 201
rect 67676 257 67732 266
rect 67676 192 67732 201
rect 68300 257 68356 266
rect 68300 192 68356 201
rect 68924 257 68980 266
rect 68924 192 68980 201
rect 69548 257 69604 266
rect 69548 192 69604 201
rect 70172 257 70228 266
rect 70172 192 70228 201
rect 70796 257 70852 266
rect 70796 192 70852 201
rect 71420 257 71476 266
rect 71420 192 71476 201
rect 72044 257 72100 266
rect 72044 192 72100 201
rect 72668 257 72724 266
rect 72668 192 72724 201
rect 73292 257 73348 266
rect 73292 192 73348 201
rect 73916 257 73972 266
rect 73916 192 73972 201
rect 74540 257 74596 266
rect 74540 192 74596 201
rect 75164 257 75220 266
rect 75164 192 75220 201
rect 75788 257 75844 266
rect 75788 192 75844 201
rect 76412 257 76468 266
rect 76412 192 76468 201
rect 77036 257 77092 266
rect 77036 192 77092 201
rect 77660 257 77716 266
rect 77660 192 77716 201
rect 78284 257 78340 266
rect 78284 192 78340 201
rect 78908 257 78964 266
rect 78908 192 78964 201
rect 79532 257 79588 266
rect 79532 192 79588 201
<< via2 >>
rect 284 201 340 257
rect 908 201 964 257
rect 1532 201 1588 257
rect 2156 201 2212 257
rect 2780 201 2836 257
rect 3404 201 3460 257
rect 4028 201 4084 257
rect 4652 201 4708 257
rect 5276 201 5332 257
rect 5900 201 5956 257
rect 6524 201 6580 257
rect 7148 201 7204 257
rect 7772 201 7828 257
rect 8396 201 8452 257
rect 9020 201 9076 257
rect 9644 201 9700 257
rect 10268 201 10324 257
rect 10892 201 10948 257
rect 11516 201 11572 257
rect 12140 201 12196 257
rect 12764 201 12820 257
rect 13388 201 13444 257
rect 14012 201 14068 257
rect 14636 201 14692 257
rect 15260 201 15316 257
rect 15884 201 15940 257
rect 16508 201 16564 257
rect 17132 201 17188 257
rect 17756 201 17812 257
rect 18380 201 18436 257
rect 19004 201 19060 257
rect 19628 201 19684 257
rect 20252 201 20308 257
rect 20876 201 20932 257
rect 21500 201 21556 257
rect 22124 201 22180 257
rect 22748 201 22804 257
rect 23372 201 23428 257
rect 23996 201 24052 257
rect 24620 201 24676 257
rect 25244 201 25300 257
rect 25868 201 25924 257
rect 26492 201 26548 257
rect 27116 201 27172 257
rect 27740 201 27796 257
rect 28364 201 28420 257
rect 28988 201 29044 257
rect 29612 201 29668 257
rect 30236 201 30292 257
rect 30860 201 30916 257
rect 31484 201 31540 257
rect 32108 201 32164 257
rect 32732 201 32788 257
rect 33356 201 33412 257
rect 33980 201 34036 257
rect 34604 201 34660 257
rect 35228 201 35284 257
rect 35852 201 35908 257
rect 36476 201 36532 257
rect 37100 201 37156 257
rect 37724 201 37780 257
rect 38348 201 38404 257
rect 38972 201 39028 257
rect 39596 201 39652 257
rect 40220 201 40276 257
rect 40844 201 40900 257
rect 41468 201 41524 257
rect 42092 201 42148 257
rect 42716 201 42772 257
rect 43340 201 43396 257
rect 43964 201 44020 257
rect 44588 201 44644 257
rect 45212 201 45268 257
rect 45836 201 45892 257
rect 46460 201 46516 257
rect 47084 201 47140 257
rect 47708 201 47764 257
rect 48332 201 48388 257
rect 48956 201 49012 257
rect 49580 201 49636 257
rect 50204 201 50260 257
rect 50828 201 50884 257
rect 51452 201 51508 257
rect 52076 201 52132 257
rect 52700 201 52756 257
rect 53324 201 53380 257
rect 53948 201 54004 257
rect 54572 201 54628 257
rect 55196 201 55252 257
rect 55820 201 55876 257
rect 56444 201 56500 257
rect 57068 201 57124 257
rect 57692 201 57748 257
rect 58316 201 58372 257
rect 58940 201 58996 257
rect 59564 201 59620 257
rect 60188 201 60244 257
rect 60812 201 60868 257
rect 61436 201 61492 257
rect 62060 201 62116 257
rect 62684 201 62740 257
rect 63308 201 63364 257
rect 63932 201 63988 257
rect 64556 201 64612 257
rect 65180 201 65236 257
rect 65804 201 65860 257
rect 66428 201 66484 257
rect 67052 201 67108 257
rect 67676 201 67732 257
rect 68300 201 68356 257
rect 68924 201 68980 257
rect 69548 201 69604 257
rect 70172 201 70228 257
rect 70796 201 70852 257
rect 71420 201 71476 257
rect 72044 201 72100 257
rect 72668 201 72724 257
rect 73292 201 73348 257
rect 73916 201 73972 257
rect 74540 201 74596 257
rect 75164 201 75220 257
rect 75788 201 75844 257
rect 76412 201 76468 257
rect 77036 201 77092 257
rect 77660 201 77716 257
rect 78284 201 78340 257
rect 78908 201 78964 257
rect 79532 201 79588 257
<< metal3 >>
rect 263 257 361 278
rect 263 201 284 257
rect 340 201 361 257
rect 263 180 361 201
rect 887 257 985 278
rect 887 201 908 257
rect 964 201 985 257
rect 887 180 985 201
rect 1511 257 1609 278
rect 1511 201 1532 257
rect 1588 201 1609 257
rect 1511 180 1609 201
rect 2135 257 2233 278
rect 2135 201 2156 257
rect 2212 201 2233 257
rect 2135 180 2233 201
rect 2759 257 2857 278
rect 2759 201 2780 257
rect 2836 201 2857 257
rect 2759 180 2857 201
rect 3383 257 3481 278
rect 3383 201 3404 257
rect 3460 201 3481 257
rect 3383 180 3481 201
rect 4007 257 4105 278
rect 4007 201 4028 257
rect 4084 201 4105 257
rect 4007 180 4105 201
rect 4631 257 4729 278
rect 4631 201 4652 257
rect 4708 201 4729 257
rect 4631 180 4729 201
rect 5255 257 5353 278
rect 5255 201 5276 257
rect 5332 201 5353 257
rect 5255 180 5353 201
rect 5879 257 5977 278
rect 5879 201 5900 257
rect 5956 201 5977 257
rect 5879 180 5977 201
rect 6503 257 6601 278
rect 6503 201 6524 257
rect 6580 201 6601 257
rect 6503 180 6601 201
rect 7127 257 7225 278
rect 7127 201 7148 257
rect 7204 201 7225 257
rect 7127 180 7225 201
rect 7751 257 7849 278
rect 7751 201 7772 257
rect 7828 201 7849 257
rect 7751 180 7849 201
rect 8375 257 8473 278
rect 8375 201 8396 257
rect 8452 201 8473 257
rect 8375 180 8473 201
rect 8999 257 9097 278
rect 8999 201 9020 257
rect 9076 201 9097 257
rect 8999 180 9097 201
rect 9623 257 9721 278
rect 9623 201 9644 257
rect 9700 201 9721 257
rect 9623 180 9721 201
rect 10247 257 10345 278
rect 10247 201 10268 257
rect 10324 201 10345 257
rect 10247 180 10345 201
rect 10871 257 10969 278
rect 10871 201 10892 257
rect 10948 201 10969 257
rect 10871 180 10969 201
rect 11495 257 11593 278
rect 11495 201 11516 257
rect 11572 201 11593 257
rect 11495 180 11593 201
rect 12119 257 12217 278
rect 12119 201 12140 257
rect 12196 201 12217 257
rect 12119 180 12217 201
rect 12743 257 12841 278
rect 12743 201 12764 257
rect 12820 201 12841 257
rect 12743 180 12841 201
rect 13367 257 13465 278
rect 13367 201 13388 257
rect 13444 201 13465 257
rect 13367 180 13465 201
rect 13991 257 14089 278
rect 13991 201 14012 257
rect 14068 201 14089 257
rect 13991 180 14089 201
rect 14615 257 14713 278
rect 14615 201 14636 257
rect 14692 201 14713 257
rect 14615 180 14713 201
rect 15239 257 15337 278
rect 15239 201 15260 257
rect 15316 201 15337 257
rect 15239 180 15337 201
rect 15863 257 15961 278
rect 15863 201 15884 257
rect 15940 201 15961 257
rect 15863 180 15961 201
rect 16487 257 16585 278
rect 16487 201 16508 257
rect 16564 201 16585 257
rect 16487 180 16585 201
rect 17111 257 17209 278
rect 17111 201 17132 257
rect 17188 201 17209 257
rect 17111 180 17209 201
rect 17735 257 17833 278
rect 17735 201 17756 257
rect 17812 201 17833 257
rect 17735 180 17833 201
rect 18359 257 18457 278
rect 18359 201 18380 257
rect 18436 201 18457 257
rect 18359 180 18457 201
rect 18983 257 19081 278
rect 18983 201 19004 257
rect 19060 201 19081 257
rect 18983 180 19081 201
rect 19607 257 19705 278
rect 19607 201 19628 257
rect 19684 201 19705 257
rect 19607 180 19705 201
rect 20231 257 20329 278
rect 20231 201 20252 257
rect 20308 201 20329 257
rect 20231 180 20329 201
rect 20855 257 20953 278
rect 20855 201 20876 257
rect 20932 201 20953 257
rect 20855 180 20953 201
rect 21479 257 21577 278
rect 21479 201 21500 257
rect 21556 201 21577 257
rect 21479 180 21577 201
rect 22103 257 22201 278
rect 22103 201 22124 257
rect 22180 201 22201 257
rect 22103 180 22201 201
rect 22727 257 22825 278
rect 22727 201 22748 257
rect 22804 201 22825 257
rect 22727 180 22825 201
rect 23351 257 23449 278
rect 23351 201 23372 257
rect 23428 201 23449 257
rect 23351 180 23449 201
rect 23975 257 24073 278
rect 23975 201 23996 257
rect 24052 201 24073 257
rect 23975 180 24073 201
rect 24599 257 24697 278
rect 24599 201 24620 257
rect 24676 201 24697 257
rect 24599 180 24697 201
rect 25223 257 25321 278
rect 25223 201 25244 257
rect 25300 201 25321 257
rect 25223 180 25321 201
rect 25847 257 25945 278
rect 25847 201 25868 257
rect 25924 201 25945 257
rect 25847 180 25945 201
rect 26471 257 26569 278
rect 26471 201 26492 257
rect 26548 201 26569 257
rect 26471 180 26569 201
rect 27095 257 27193 278
rect 27095 201 27116 257
rect 27172 201 27193 257
rect 27095 180 27193 201
rect 27719 257 27817 278
rect 27719 201 27740 257
rect 27796 201 27817 257
rect 27719 180 27817 201
rect 28343 257 28441 278
rect 28343 201 28364 257
rect 28420 201 28441 257
rect 28343 180 28441 201
rect 28967 257 29065 278
rect 28967 201 28988 257
rect 29044 201 29065 257
rect 28967 180 29065 201
rect 29591 257 29689 278
rect 29591 201 29612 257
rect 29668 201 29689 257
rect 29591 180 29689 201
rect 30215 257 30313 278
rect 30215 201 30236 257
rect 30292 201 30313 257
rect 30215 180 30313 201
rect 30839 257 30937 278
rect 30839 201 30860 257
rect 30916 201 30937 257
rect 30839 180 30937 201
rect 31463 257 31561 278
rect 31463 201 31484 257
rect 31540 201 31561 257
rect 31463 180 31561 201
rect 32087 257 32185 278
rect 32087 201 32108 257
rect 32164 201 32185 257
rect 32087 180 32185 201
rect 32711 257 32809 278
rect 32711 201 32732 257
rect 32788 201 32809 257
rect 32711 180 32809 201
rect 33335 257 33433 278
rect 33335 201 33356 257
rect 33412 201 33433 257
rect 33335 180 33433 201
rect 33959 257 34057 278
rect 33959 201 33980 257
rect 34036 201 34057 257
rect 33959 180 34057 201
rect 34583 257 34681 278
rect 34583 201 34604 257
rect 34660 201 34681 257
rect 34583 180 34681 201
rect 35207 257 35305 278
rect 35207 201 35228 257
rect 35284 201 35305 257
rect 35207 180 35305 201
rect 35831 257 35929 278
rect 35831 201 35852 257
rect 35908 201 35929 257
rect 35831 180 35929 201
rect 36455 257 36553 278
rect 36455 201 36476 257
rect 36532 201 36553 257
rect 36455 180 36553 201
rect 37079 257 37177 278
rect 37079 201 37100 257
rect 37156 201 37177 257
rect 37079 180 37177 201
rect 37703 257 37801 278
rect 37703 201 37724 257
rect 37780 201 37801 257
rect 37703 180 37801 201
rect 38327 257 38425 278
rect 38327 201 38348 257
rect 38404 201 38425 257
rect 38327 180 38425 201
rect 38951 257 39049 278
rect 38951 201 38972 257
rect 39028 201 39049 257
rect 38951 180 39049 201
rect 39575 257 39673 278
rect 39575 201 39596 257
rect 39652 201 39673 257
rect 39575 180 39673 201
rect 40199 257 40297 278
rect 40199 201 40220 257
rect 40276 201 40297 257
rect 40199 180 40297 201
rect 40823 257 40921 278
rect 40823 201 40844 257
rect 40900 201 40921 257
rect 40823 180 40921 201
rect 41447 257 41545 278
rect 41447 201 41468 257
rect 41524 201 41545 257
rect 41447 180 41545 201
rect 42071 257 42169 278
rect 42071 201 42092 257
rect 42148 201 42169 257
rect 42071 180 42169 201
rect 42695 257 42793 278
rect 42695 201 42716 257
rect 42772 201 42793 257
rect 42695 180 42793 201
rect 43319 257 43417 278
rect 43319 201 43340 257
rect 43396 201 43417 257
rect 43319 180 43417 201
rect 43943 257 44041 278
rect 43943 201 43964 257
rect 44020 201 44041 257
rect 43943 180 44041 201
rect 44567 257 44665 278
rect 44567 201 44588 257
rect 44644 201 44665 257
rect 44567 180 44665 201
rect 45191 257 45289 278
rect 45191 201 45212 257
rect 45268 201 45289 257
rect 45191 180 45289 201
rect 45815 257 45913 278
rect 45815 201 45836 257
rect 45892 201 45913 257
rect 45815 180 45913 201
rect 46439 257 46537 278
rect 46439 201 46460 257
rect 46516 201 46537 257
rect 46439 180 46537 201
rect 47063 257 47161 278
rect 47063 201 47084 257
rect 47140 201 47161 257
rect 47063 180 47161 201
rect 47687 257 47785 278
rect 47687 201 47708 257
rect 47764 201 47785 257
rect 47687 180 47785 201
rect 48311 257 48409 278
rect 48311 201 48332 257
rect 48388 201 48409 257
rect 48311 180 48409 201
rect 48935 257 49033 278
rect 48935 201 48956 257
rect 49012 201 49033 257
rect 48935 180 49033 201
rect 49559 257 49657 278
rect 49559 201 49580 257
rect 49636 201 49657 257
rect 49559 180 49657 201
rect 50183 257 50281 278
rect 50183 201 50204 257
rect 50260 201 50281 257
rect 50183 180 50281 201
rect 50807 257 50905 278
rect 50807 201 50828 257
rect 50884 201 50905 257
rect 50807 180 50905 201
rect 51431 257 51529 278
rect 51431 201 51452 257
rect 51508 201 51529 257
rect 51431 180 51529 201
rect 52055 257 52153 278
rect 52055 201 52076 257
rect 52132 201 52153 257
rect 52055 180 52153 201
rect 52679 257 52777 278
rect 52679 201 52700 257
rect 52756 201 52777 257
rect 52679 180 52777 201
rect 53303 257 53401 278
rect 53303 201 53324 257
rect 53380 201 53401 257
rect 53303 180 53401 201
rect 53927 257 54025 278
rect 53927 201 53948 257
rect 54004 201 54025 257
rect 53927 180 54025 201
rect 54551 257 54649 278
rect 54551 201 54572 257
rect 54628 201 54649 257
rect 54551 180 54649 201
rect 55175 257 55273 278
rect 55175 201 55196 257
rect 55252 201 55273 257
rect 55175 180 55273 201
rect 55799 257 55897 278
rect 55799 201 55820 257
rect 55876 201 55897 257
rect 55799 180 55897 201
rect 56423 257 56521 278
rect 56423 201 56444 257
rect 56500 201 56521 257
rect 56423 180 56521 201
rect 57047 257 57145 278
rect 57047 201 57068 257
rect 57124 201 57145 257
rect 57047 180 57145 201
rect 57671 257 57769 278
rect 57671 201 57692 257
rect 57748 201 57769 257
rect 57671 180 57769 201
rect 58295 257 58393 278
rect 58295 201 58316 257
rect 58372 201 58393 257
rect 58295 180 58393 201
rect 58919 257 59017 278
rect 58919 201 58940 257
rect 58996 201 59017 257
rect 58919 180 59017 201
rect 59543 257 59641 278
rect 59543 201 59564 257
rect 59620 201 59641 257
rect 59543 180 59641 201
rect 60167 257 60265 278
rect 60167 201 60188 257
rect 60244 201 60265 257
rect 60167 180 60265 201
rect 60791 257 60889 278
rect 60791 201 60812 257
rect 60868 201 60889 257
rect 60791 180 60889 201
rect 61415 257 61513 278
rect 61415 201 61436 257
rect 61492 201 61513 257
rect 61415 180 61513 201
rect 62039 257 62137 278
rect 62039 201 62060 257
rect 62116 201 62137 257
rect 62039 180 62137 201
rect 62663 257 62761 278
rect 62663 201 62684 257
rect 62740 201 62761 257
rect 62663 180 62761 201
rect 63287 257 63385 278
rect 63287 201 63308 257
rect 63364 201 63385 257
rect 63287 180 63385 201
rect 63911 257 64009 278
rect 63911 201 63932 257
rect 63988 201 64009 257
rect 63911 180 64009 201
rect 64535 257 64633 278
rect 64535 201 64556 257
rect 64612 201 64633 257
rect 64535 180 64633 201
rect 65159 257 65257 278
rect 65159 201 65180 257
rect 65236 201 65257 257
rect 65159 180 65257 201
rect 65783 257 65881 278
rect 65783 201 65804 257
rect 65860 201 65881 257
rect 65783 180 65881 201
rect 66407 257 66505 278
rect 66407 201 66428 257
rect 66484 201 66505 257
rect 66407 180 66505 201
rect 67031 257 67129 278
rect 67031 201 67052 257
rect 67108 201 67129 257
rect 67031 180 67129 201
rect 67655 257 67753 278
rect 67655 201 67676 257
rect 67732 201 67753 257
rect 67655 180 67753 201
rect 68279 257 68377 278
rect 68279 201 68300 257
rect 68356 201 68377 257
rect 68279 180 68377 201
rect 68903 257 69001 278
rect 68903 201 68924 257
rect 68980 201 69001 257
rect 68903 180 69001 201
rect 69527 257 69625 278
rect 69527 201 69548 257
rect 69604 201 69625 257
rect 69527 180 69625 201
rect 70151 257 70249 278
rect 70151 201 70172 257
rect 70228 201 70249 257
rect 70151 180 70249 201
rect 70775 257 70873 278
rect 70775 201 70796 257
rect 70852 201 70873 257
rect 70775 180 70873 201
rect 71399 257 71497 278
rect 71399 201 71420 257
rect 71476 201 71497 257
rect 71399 180 71497 201
rect 72023 257 72121 278
rect 72023 201 72044 257
rect 72100 201 72121 257
rect 72023 180 72121 201
rect 72647 257 72745 278
rect 72647 201 72668 257
rect 72724 201 72745 257
rect 72647 180 72745 201
rect 73271 257 73369 278
rect 73271 201 73292 257
rect 73348 201 73369 257
rect 73271 180 73369 201
rect 73895 257 73993 278
rect 73895 201 73916 257
rect 73972 201 73993 257
rect 73895 180 73993 201
rect 74519 257 74617 278
rect 74519 201 74540 257
rect 74596 201 74617 257
rect 74519 180 74617 201
rect 75143 257 75241 278
rect 75143 201 75164 257
rect 75220 201 75241 257
rect 75143 180 75241 201
rect 75767 257 75865 278
rect 75767 201 75788 257
rect 75844 201 75865 257
rect 75767 180 75865 201
rect 76391 257 76489 278
rect 76391 201 76412 257
rect 76468 201 76489 257
rect 76391 180 76489 201
rect 77015 257 77113 278
rect 77015 201 77036 257
rect 77092 201 77113 257
rect 77015 180 77113 201
rect 77639 257 77737 278
rect 77639 201 77660 257
rect 77716 201 77737 257
rect 77639 180 77737 201
rect 78263 257 78361 278
rect 78263 201 78284 257
rect 78340 201 78361 257
rect 78263 180 78361 201
rect 78887 257 78985 278
rect 78887 201 78908 257
rect 78964 201 78985 257
rect 78887 180 78985 201
rect 79511 257 79609 278
rect 79511 201 79532 257
rect 79588 201 79609 257
rect 79511 180 79609 201
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_0
timestamp 1676037725
transform -1 0 19968 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_1
timestamp 1676037725
transform 1 0 18720 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_2
timestamp 1676037725
transform -1 0 18720 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_3
timestamp 1676037725
transform 1 0 17472 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_4
timestamp 1676037725
transform -1 0 17472 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_5
timestamp 1676037725
transform 1 0 16224 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_6
timestamp 1676037725
transform -1 0 16224 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_7
timestamp 1676037725
transform 1 0 14976 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_8
timestamp 1676037725
transform -1 0 14976 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_9
timestamp 1676037725
transform 1 0 13728 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_10
timestamp 1676037725
transform -1 0 13728 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_11
timestamp 1676037725
transform 1 0 12480 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_12
timestamp 1676037725
transform -1 0 12480 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_13
timestamp 1676037725
transform 1 0 11232 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_14
timestamp 1676037725
transform -1 0 11232 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_15
timestamp 1676037725
transform 1 0 9984 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_16
timestamp 1676037725
transform -1 0 9984 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_17
timestamp 1676037725
transform 1 0 8736 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_18
timestamp 1676037725
transform -1 0 8736 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_19
timestamp 1676037725
transform 1 0 7488 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_20
timestamp 1676037725
transform -1 0 7488 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_21
timestamp 1676037725
transform 1 0 6240 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_22
timestamp 1676037725
transform -1 0 6240 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_23
timestamp 1676037725
transform 1 0 4992 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_24
timestamp 1676037725
transform -1 0 4992 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_25
timestamp 1676037725
transform 1 0 3744 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_26
timestamp 1676037725
transform -1 0 3744 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_27
timestamp 1676037725
transform 1 0 2496 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_28
timestamp 1676037725
transform -1 0 2496 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_29
timestamp 1676037725
transform 1 0 1248 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_30
timestamp 1676037725
transform -1 0 1248 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_31
timestamp 1676037725
transform 1 0 0 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_32
timestamp 1676037725
transform -1 0 39936 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_33
timestamp 1676037725
transform 1 0 38688 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_34
timestamp 1676037725
transform -1 0 38688 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_35
timestamp 1676037725
transform 1 0 37440 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_36
timestamp 1676037725
transform -1 0 37440 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_37
timestamp 1676037725
transform 1 0 36192 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_38
timestamp 1676037725
transform -1 0 36192 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_39
timestamp 1676037725
transform 1 0 34944 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_40
timestamp 1676037725
transform -1 0 34944 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_41
timestamp 1676037725
transform 1 0 33696 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_42
timestamp 1676037725
transform -1 0 33696 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_43
timestamp 1676037725
transform 1 0 32448 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_44
timestamp 1676037725
transform -1 0 32448 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_45
timestamp 1676037725
transform 1 0 31200 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_46
timestamp 1676037725
transform -1 0 31200 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_47
timestamp 1676037725
transform 1 0 29952 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_48
timestamp 1676037725
transform -1 0 29952 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_49
timestamp 1676037725
transform 1 0 28704 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_50
timestamp 1676037725
transform -1 0 28704 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_51
timestamp 1676037725
transform 1 0 27456 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_52
timestamp 1676037725
transform -1 0 27456 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_53
timestamp 1676037725
transform 1 0 26208 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_54
timestamp 1676037725
transform -1 0 26208 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_55
timestamp 1676037725
transform 1 0 24960 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_56
timestamp 1676037725
transform -1 0 24960 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_57
timestamp 1676037725
transform 1 0 23712 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_58
timestamp 1676037725
transform -1 0 23712 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_59
timestamp 1676037725
transform 1 0 22464 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_60
timestamp 1676037725
transform -1 0 22464 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_61
timestamp 1676037725
transform 1 0 21216 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_62
timestamp 1676037725
transform -1 0 21216 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_63
timestamp 1676037725
transform 1 0 19968 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_64
timestamp 1676037725
transform -1 0 59904 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_65
timestamp 1676037725
transform 1 0 58656 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_66
timestamp 1676037725
transform -1 0 58656 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_67
timestamp 1676037725
transform 1 0 57408 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_68
timestamp 1676037725
transform -1 0 57408 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_69
timestamp 1676037725
transform 1 0 56160 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_70
timestamp 1676037725
transform -1 0 56160 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_71
timestamp 1676037725
transform 1 0 54912 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_72
timestamp 1676037725
transform -1 0 54912 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_73
timestamp 1676037725
transform 1 0 53664 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_74
timestamp 1676037725
transform -1 0 53664 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_75
timestamp 1676037725
transform 1 0 52416 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_76
timestamp 1676037725
transform -1 0 52416 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_77
timestamp 1676037725
transform 1 0 51168 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_78
timestamp 1676037725
transform -1 0 51168 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_79
timestamp 1676037725
transform 1 0 49920 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_80
timestamp 1676037725
transform -1 0 49920 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_81
timestamp 1676037725
transform 1 0 48672 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_82
timestamp 1676037725
transform -1 0 48672 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_83
timestamp 1676037725
transform 1 0 47424 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_84
timestamp 1676037725
transform -1 0 47424 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_85
timestamp 1676037725
transform 1 0 46176 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_86
timestamp 1676037725
transform -1 0 46176 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_87
timestamp 1676037725
transform 1 0 44928 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_88
timestamp 1676037725
transform -1 0 44928 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_89
timestamp 1676037725
transform 1 0 43680 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_90
timestamp 1676037725
transform -1 0 43680 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_91
timestamp 1676037725
transform 1 0 42432 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_92
timestamp 1676037725
transform -1 0 42432 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_93
timestamp 1676037725
transform 1 0 41184 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_94
timestamp 1676037725
transform -1 0 41184 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_95
timestamp 1676037725
transform 1 0 39936 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_96
timestamp 1676037725
transform -1 0 79872 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_97
timestamp 1676037725
transform 1 0 78624 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_98
timestamp 1676037725
transform -1 0 78624 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_99
timestamp 1676037725
transform 1 0 77376 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_100
timestamp 1676037725
transform -1 0 77376 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_101
timestamp 1676037725
transform 1 0 76128 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_102
timestamp 1676037725
transform -1 0 76128 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_103
timestamp 1676037725
transform 1 0 74880 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_104
timestamp 1676037725
transform -1 0 74880 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_105
timestamp 1676037725
transform 1 0 73632 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_106
timestamp 1676037725
transform -1 0 73632 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_107
timestamp 1676037725
transform 1 0 72384 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_108
timestamp 1676037725
transform -1 0 72384 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_109
timestamp 1676037725
transform 1 0 71136 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_110
timestamp 1676037725
transform -1 0 71136 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_111
timestamp 1676037725
transform 1 0 69888 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_112
timestamp 1676037725
transform -1 0 69888 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_113
timestamp 1676037725
transform 1 0 68640 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_114
timestamp 1676037725
transform -1 0 68640 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_115
timestamp 1676037725
transform 1 0 67392 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_116
timestamp 1676037725
transform -1 0 67392 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_117
timestamp 1676037725
transform 1 0 66144 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_118
timestamp 1676037725
transform -1 0 66144 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_119
timestamp 1676037725
transform 1 0 64896 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_120
timestamp 1676037725
transform -1 0 64896 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_121
timestamp 1676037725
transform 1 0 63648 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_122
timestamp 1676037725
transform -1 0 63648 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_123
timestamp 1676037725
transform 1 0 62400 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_124
timestamp 1676037725
transform -1 0 62400 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_125
timestamp 1676037725
transform 1 0 61152 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_126
timestamp 1676037725
transform -1 0 61152 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_127
timestamp 1676037725
transform 1 0 59904 0 1 0
box 0 0 624 474
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1676037725
transform 1 0 19623 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1676037725
transform 1 0 18999 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1676037725
transform 1 0 18375 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1676037725
transform 1 0 17751 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1676037725
transform 1 0 17127 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1676037725
transform 1 0 16503 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1676037725
transform 1 0 15879 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1676037725
transform 1 0 15255 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1676037725
transform 1 0 14631 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1676037725
transform 1 0 14007 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1676037725
transform 1 0 13383 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1676037725
transform 1 0 12759 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1676037725
transform 1 0 12135 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1676037725
transform 1 0 11511 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1676037725
transform 1 0 10887 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1676037725
transform 1 0 10263 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1676037725
transform 1 0 9639 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1676037725
transform 1 0 9015 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1676037725
transform 1 0 8391 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1676037725
transform 1 0 7767 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1676037725
transform 1 0 7143 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1676037725
transform 1 0 6519 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1676037725
transform 1 0 5895 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1676037725
transform 1 0 5271 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1676037725
transform 1 0 4647 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1676037725
transform 1 0 4023 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1676037725
transform 1 0 3399 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1676037725
transform 1 0 2775 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1676037725
transform 1 0 2151 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1676037725
transform 1 0 1527 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1676037725
transform 1 0 903 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1676037725
transform 1 0 279 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1676037725
transform 1 0 39591 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1676037725
transform 1 0 38967 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1676037725
transform 1 0 38343 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1676037725
transform 1 0 37719 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1676037725
transform 1 0 37095 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1676037725
transform 1 0 36471 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1676037725
transform 1 0 35847 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1676037725
transform 1 0 35223 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1676037725
transform 1 0 34599 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1676037725
transform 1 0 33975 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1676037725
transform 1 0 33351 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1676037725
transform 1 0 32727 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1676037725
transform 1 0 32103 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1676037725
transform 1 0 31479 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1676037725
transform 1 0 30855 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1676037725
transform 1 0 30231 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1676037725
transform 1 0 29607 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1676037725
transform 1 0 28983 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1676037725
transform 1 0 28359 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1676037725
transform 1 0 27735 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1676037725
transform 1 0 27111 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1676037725
transform 1 0 26487 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1676037725
transform 1 0 25863 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1676037725
transform 1 0 25239 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1676037725
transform 1 0 24615 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1676037725
transform 1 0 23991 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1676037725
transform 1 0 23367 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1676037725
transform 1 0 22743 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1676037725
transform 1 0 22119 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1676037725
transform 1 0 21495 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1676037725
transform 1 0 20871 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1676037725
transform 1 0 20247 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1676037725
transform 1 0 59559 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1676037725
transform 1 0 58935 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1676037725
transform 1 0 58311 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1676037725
transform 1 0 57687 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1676037725
transform 1 0 57063 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1676037725
transform 1 0 56439 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1676037725
transform 1 0 55815 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1676037725
transform 1 0 55191 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_72
timestamp 1676037725
transform 1 0 54567 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_73
timestamp 1676037725
transform 1 0 53943 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_74
timestamp 1676037725
transform 1 0 53319 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_75
timestamp 1676037725
transform 1 0 52695 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_76
timestamp 1676037725
transform 1 0 52071 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_77
timestamp 1676037725
transform 1 0 51447 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_78
timestamp 1676037725
transform 1 0 50823 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_79
timestamp 1676037725
transform 1 0 50199 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_80
timestamp 1676037725
transform 1 0 49575 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_81
timestamp 1676037725
transform 1 0 48951 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_82
timestamp 1676037725
transform 1 0 48327 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_83
timestamp 1676037725
transform 1 0 47703 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_84
timestamp 1676037725
transform 1 0 47079 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_85
timestamp 1676037725
transform 1 0 46455 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_86
timestamp 1676037725
transform 1 0 45831 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_87
timestamp 1676037725
transform 1 0 45207 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_88
timestamp 1676037725
transform 1 0 44583 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_89
timestamp 1676037725
transform 1 0 43959 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_90
timestamp 1676037725
transform 1 0 43335 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_91
timestamp 1676037725
transform 1 0 42711 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_92
timestamp 1676037725
transform 1 0 42087 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_93
timestamp 1676037725
transform 1 0 41463 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_94
timestamp 1676037725
transform 1 0 40839 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_95
timestamp 1676037725
transform 1 0 40215 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_96
timestamp 1676037725
transform 1 0 79527 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_97
timestamp 1676037725
transform 1 0 78903 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_98
timestamp 1676037725
transform 1 0 78279 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_99
timestamp 1676037725
transform 1 0 77655 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_100
timestamp 1676037725
transform 1 0 77031 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_101
timestamp 1676037725
transform 1 0 76407 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_102
timestamp 1676037725
transform 1 0 75783 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_103
timestamp 1676037725
transform 1 0 75159 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_104
timestamp 1676037725
transform 1 0 74535 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_105
timestamp 1676037725
transform 1 0 73911 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_106
timestamp 1676037725
transform 1 0 73287 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_107
timestamp 1676037725
transform 1 0 72663 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_108
timestamp 1676037725
transform 1 0 72039 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_109
timestamp 1676037725
transform 1 0 71415 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_110
timestamp 1676037725
transform 1 0 70791 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_111
timestamp 1676037725
transform 1 0 70167 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_112
timestamp 1676037725
transform 1 0 69543 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_113
timestamp 1676037725
transform 1 0 68919 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_114
timestamp 1676037725
transform 1 0 68295 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_115
timestamp 1676037725
transform 1 0 67671 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_116
timestamp 1676037725
transform 1 0 67047 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_117
timestamp 1676037725
transform 1 0 66423 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_118
timestamp 1676037725
transform 1 0 65799 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_119
timestamp 1676037725
transform 1 0 65175 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_120
timestamp 1676037725
transform 1 0 64551 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_121
timestamp 1676037725
transform 1 0 63927 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_122
timestamp 1676037725
transform 1 0 63303 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_123
timestamp 1676037725
transform 1 0 62679 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_124
timestamp 1676037725
transform 1 0 62055 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_125
timestamp 1676037725
transform 1 0 61431 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_126
timestamp 1676037725
transform 1 0 60807 0 1 192
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_127
timestamp 1676037725
transform 1 0 60183 0 1 192
box 0 0 1 1
<< labels >>
rlabel metal3 s 29591 180 29689 278 4 vdd
rlabel metal3 s 20231 180 20329 278 4 vdd
rlabel metal3 s 20855 180 20953 278 4 vdd
rlabel metal3 s 14615 180 14713 278 4 vdd
rlabel metal3 s 6503 180 6601 278 4 vdd
rlabel metal3 s 5879 180 5977 278 4 vdd
rlabel metal3 s 32087 180 32185 278 4 vdd
rlabel metal3 s 25223 180 25321 278 4 vdd
rlabel metal3 s 15863 180 15961 278 4 vdd
rlabel metal3 s 15239 180 15337 278 4 vdd
rlabel metal3 s 17111 180 17209 278 4 vdd
rlabel metal3 s 2759 180 2857 278 4 vdd
rlabel metal3 s 19607 180 19705 278 4 vdd
rlabel metal3 s 26471 180 26569 278 4 vdd
rlabel metal3 s 38951 180 39049 278 4 vdd
rlabel metal3 s 22103 180 22201 278 4 vdd
rlabel metal3 s 7751 180 7849 278 4 vdd
rlabel metal3 s 31463 180 31561 278 4 vdd
rlabel metal3 s 21479 180 21577 278 4 vdd
rlabel metal3 s 10247 180 10345 278 4 vdd
rlabel metal3 s 33335 180 33433 278 4 vdd
rlabel metal3 s 4007 180 4105 278 4 vdd
rlabel metal3 s 8999 180 9097 278 4 vdd
rlabel metal3 s 24599 180 24697 278 4 vdd
rlabel metal3 s 38327 180 38425 278 4 vdd
rlabel metal3 s 39575 180 39673 278 4 vdd
rlabel metal3 s 33959 180 34057 278 4 vdd
rlabel metal3 s 2135 180 2233 278 4 vdd
rlabel metal3 s 25847 180 25945 278 4 vdd
rlabel metal3 s 28967 180 29065 278 4 vdd
rlabel metal3 s 30839 180 30937 278 4 vdd
rlabel metal3 s 27719 180 27817 278 4 vdd
rlabel metal3 s 37079 180 37177 278 4 vdd
rlabel metal3 s 7127 180 7225 278 4 vdd
rlabel metal3 s 18359 180 18457 278 4 vdd
rlabel metal3 s 12743 180 12841 278 4 vdd
rlabel metal3 s 1511 180 1609 278 4 vdd
rlabel metal3 s 35207 180 35305 278 4 vdd
rlabel metal3 s 30215 180 30313 278 4 vdd
rlabel metal3 s 23351 180 23449 278 4 vdd
rlabel metal3 s 9623 180 9721 278 4 vdd
rlabel metal3 s 13991 180 14089 278 4 vdd
rlabel metal3 s 887 180 985 278 4 vdd
rlabel metal3 s 22727 180 22825 278 4 vdd
rlabel metal3 s 36455 180 36553 278 4 vdd
rlabel metal3 s 3383 180 3481 278 4 vdd
rlabel metal3 s 8375 180 8473 278 4 vdd
rlabel metal3 s 35831 180 35929 278 4 vdd
rlabel metal3 s 17735 180 17833 278 4 vdd
rlabel metal3 s 11495 180 11593 278 4 vdd
rlabel metal3 s 263 180 361 278 4 vdd
rlabel metal3 s 28343 180 28441 278 4 vdd
rlabel metal3 s 37703 180 37801 278 4 vdd
rlabel metal3 s 23975 180 24073 278 4 vdd
rlabel metal3 s 12119 180 12217 278 4 vdd
rlabel metal3 s 13367 180 13465 278 4 vdd
rlabel metal3 s 34583 180 34681 278 4 vdd
rlabel metal3 s 27095 180 27193 278 4 vdd
rlabel metal3 s 4631 180 4729 278 4 vdd
rlabel metal3 s 16487 180 16585 278 4 vdd
rlabel metal3 s 10871 180 10969 278 4 vdd
rlabel metal3 s 5255 180 5353 278 4 vdd
rlabel metal3 s 18983 180 19081 278 4 vdd
rlabel metal3 s 32711 180 32809 278 4 vdd
rlabel metal3 s 71399 180 71497 278 4 vdd
rlabel metal3 s 74519 180 74617 278 4 vdd
rlabel metal3 s 50183 180 50281 278 4 vdd
rlabel metal3 s 61415 180 61513 278 4 vdd
rlabel metal3 s 75767 180 75865 278 4 vdd
rlabel metal3 s 52679 180 52777 278 4 vdd
rlabel metal3 s 58295 180 58393 278 4 vdd
rlabel metal3 s 60791 180 60889 278 4 vdd
rlabel metal3 s 73271 180 73369 278 4 vdd
rlabel metal3 s 75143 180 75241 278 4 vdd
rlabel metal3 s 58919 180 59017 278 4 vdd
rlabel metal3 s 78263 180 78361 278 4 vdd
rlabel metal3 s 48311 180 48409 278 4 vdd
rlabel metal3 s 47687 180 47785 278 4 vdd
rlabel metal3 s 65783 180 65881 278 4 vdd
rlabel metal3 s 73895 180 73993 278 4 vdd
rlabel metal3 s 77639 180 77737 278 4 vdd
rlabel metal3 s 66407 180 66505 278 4 vdd
rlabel metal3 s 53303 180 53401 278 4 vdd
rlabel metal3 s 51431 180 51529 278 4 vdd
rlabel metal3 s 77015 180 77113 278 4 vdd
rlabel metal3 s 45815 180 45913 278 4 vdd
rlabel metal3 s 40199 180 40297 278 4 vdd
rlabel metal3 s 57671 180 57769 278 4 vdd
rlabel metal3 s 72647 180 72745 278 4 vdd
rlabel metal3 s 67031 180 67129 278 4 vdd
rlabel metal3 s 46439 180 46537 278 4 vdd
rlabel metal3 s 76391 180 76489 278 4 vdd
rlabel metal3 s 52055 180 52153 278 4 vdd
rlabel metal3 s 67655 180 67753 278 4 vdd
rlabel metal3 s 72023 180 72121 278 4 vdd
rlabel metal3 s 60167 180 60265 278 4 vdd
rlabel metal3 s 70775 180 70873 278 4 vdd
rlabel metal3 s 78887 180 78985 278 4 vdd
rlabel metal3 s 54551 180 54649 278 4 vdd
rlabel metal3 s 43943 180 44041 278 4 vdd
rlabel metal3 s 64535 180 64633 278 4 vdd
rlabel metal3 s 49559 180 49657 278 4 vdd
rlabel metal3 s 43319 180 43417 278 4 vdd
rlabel metal3 s 50807 180 50905 278 4 vdd
rlabel metal3 s 47063 180 47161 278 4 vdd
rlabel metal3 s 68279 180 68377 278 4 vdd
rlabel metal3 s 41447 180 41545 278 4 vdd
rlabel metal3 s 63911 180 64009 278 4 vdd
rlabel metal3 s 79511 180 79609 278 4 vdd
rlabel metal3 s 65159 180 65257 278 4 vdd
rlabel metal3 s 68903 180 69001 278 4 vdd
rlabel metal3 s 55799 180 55897 278 4 vdd
rlabel metal3 s 63287 180 63385 278 4 vdd
rlabel metal3 s 59543 180 59641 278 4 vdd
rlabel metal3 s 40823 180 40921 278 4 vdd
rlabel metal3 s 57047 180 57145 278 4 vdd
rlabel metal3 s 62663 180 62761 278 4 vdd
rlabel metal3 s 45191 180 45289 278 4 vdd
rlabel metal3 s 70151 180 70249 278 4 vdd
rlabel metal3 s 42695 180 42793 278 4 vdd
rlabel metal3 s 48935 180 49033 278 4 vdd
rlabel metal3 s 53927 180 54025 278 4 vdd
rlabel metal3 s 44567 180 44665 278 4 vdd
rlabel metal3 s 56423 180 56521 278 4 vdd
rlabel metal3 s 55175 180 55273 278 4 vdd
rlabel metal3 s 42071 180 42169 278 4 vdd
rlabel metal3 s 62039 180 62137 278 4 vdd
rlabel metal3 s 69527 180 69625 278 4 vdd
rlabel metal1 s 78 0 114 395 4 bl0_0
rlabel metal1 s 150 0 186 395 4 br0_0
rlabel metal1 s 294 0 330 395 4 bl1_0
rlabel metal1 s 366 0 402 395 4 br1_0
rlabel metal1 s 1134 0 1170 395 4 bl0_1
rlabel metal1 s 1062 0 1098 395 4 br0_1
rlabel metal1 s 918 0 954 395 4 bl1_1
rlabel metal1 s 846 0 882 395 4 br1_1
rlabel metal1 s 1326 0 1362 395 4 bl0_2
rlabel metal1 s 1398 0 1434 395 4 br0_2
rlabel metal1 s 1542 0 1578 395 4 bl1_2
rlabel metal1 s 1614 0 1650 395 4 br1_2
rlabel metal1 s 2382 0 2418 395 4 bl0_3
rlabel metal1 s 2310 0 2346 395 4 br0_3
rlabel metal1 s 2166 0 2202 395 4 bl1_3
rlabel metal1 s 2094 0 2130 395 4 br1_3
rlabel metal1 s 2574 0 2610 395 4 bl0_4
rlabel metal1 s 2646 0 2682 395 4 br0_4
rlabel metal1 s 2790 0 2826 395 4 bl1_4
rlabel metal1 s 2862 0 2898 395 4 br1_4
rlabel metal1 s 3630 0 3666 395 4 bl0_5
rlabel metal1 s 3558 0 3594 395 4 br0_5
rlabel metal1 s 3414 0 3450 395 4 bl1_5
rlabel metal1 s 3342 0 3378 395 4 br1_5
rlabel metal1 s 3822 0 3858 395 4 bl0_6
rlabel metal1 s 3894 0 3930 395 4 br0_6
rlabel metal1 s 4038 0 4074 395 4 bl1_6
rlabel metal1 s 4110 0 4146 395 4 br1_6
rlabel metal1 s 4878 0 4914 395 4 bl0_7
rlabel metal1 s 4806 0 4842 395 4 br0_7
rlabel metal1 s 4662 0 4698 395 4 bl1_7
rlabel metal1 s 4590 0 4626 395 4 br1_7
rlabel metal1 s 5070 0 5106 395 4 bl0_8
rlabel metal1 s 5142 0 5178 395 4 br0_8
rlabel metal1 s 5286 0 5322 395 4 bl1_8
rlabel metal1 s 5358 0 5394 395 4 br1_8
rlabel metal1 s 6126 0 6162 395 4 bl0_9
rlabel metal1 s 6054 0 6090 395 4 br0_9
rlabel metal1 s 5910 0 5946 395 4 bl1_9
rlabel metal1 s 5838 0 5874 395 4 br1_9
rlabel metal1 s 6318 0 6354 395 4 bl0_10
rlabel metal1 s 6390 0 6426 395 4 br0_10
rlabel metal1 s 6534 0 6570 395 4 bl1_10
rlabel metal1 s 6606 0 6642 395 4 br1_10
rlabel metal1 s 7374 0 7410 395 4 bl0_11
rlabel metal1 s 7302 0 7338 395 4 br0_11
rlabel metal1 s 7158 0 7194 395 4 bl1_11
rlabel metal1 s 7086 0 7122 395 4 br1_11
rlabel metal1 s 7566 0 7602 395 4 bl0_12
rlabel metal1 s 7638 0 7674 395 4 br0_12
rlabel metal1 s 7782 0 7818 395 4 bl1_12
rlabel metal1 s 7854 0 7890 395 4 br1_12
rlabel metal1 s 8622 0 8658 395 4 bl0_13
rlabel metal1 s 8550 0 8586 395 4 br0_13
rlabel metal1 s 8406 0 8442 395 4 bl1_13
rlabel metal1 s 8334 0 8370 395 4 br1_13
rlabel metal1 s 8814 0 8850 395 4 bl0_14
rlabel metal1 s 8886 0 8922 395 4 br0_14
rlabel metal1 s 9030 0 9066 395 4 bl1_14
rlabel metal1 s 9102 0 9138 395 4 br1_14
rlabel metal1 s 9870 0 9906 395 4 bl0_15
rlabel metal1 s 9798 0 9834 395 4 br0_15
rlabel metal1 s 9654 0 9690 395 4 bl1_15
rlabel metal1 s 9582 0 9618 395 4 br1_15
rlabel metal1 s 10062 0 10098 395 4 bl0_16
rlabel metal1 s 10134 0 10170 395 4 br0_16
rlabel metal1 s 10278 0 10314 395 4 bl1_16
rlabel metal1 s 10350 0 10386 395 4 br1_16
rlabel metal1 s 11118 0 11154 395 4 bl0_17
rlabel metal1 s 11046 0 11082 395 4 br0_17
rlabel metal1 s 10902 0 10938 395 4 bl1_17
rlabel metal1 s 10830 0 10866 395 4 br1_17
rlabel metal1 s 11310 0 11346 395 4 bl0_18
rlabel metal1 s 11382 0 11418 395 4 br0_18
rlabel metal1 s 11526 0 11562 395 4 bl1_18
rlabel metal1 s 11598 0 11634 395 4 br1_18
rlabel metal1 s 12366 0 12402 395 4 bl0_19
rlabel metal1 s 12294 0 12330 395 4 br0_19
rlabel metal1 s 12150 0 12186 395 4 bl1_19
rlabel metal1 s 12078 0 12114 395 4 br1_19
rlabel metal1 s 12558 0 12594 395 4 bl0_20
rlabel metal1 s 12630 0 12666 395 4 br0_20
rlabel metal1 s 12774 0 12810 395 4 bl1_20
rlabel metal1 s 12846 0 12882 395 4 br1_20
rlabel metal1 s 13614 0 13650 395 4 bl0_21
rlabel metal1 s 13542 0 13578 395 4 br0_21
rlabel metal1 s 13398 0 13434 395 4 bl1_21
rlabel metal1 s 13326 0 13362 395 4 br1_21
rlabel metal1 s 13806 0 13842 395 4 bl0_22
rlabel metal1 s 13878 0 13914 395 4 br0_22
rlabel metal1 s 14022 0 14058 395 4 bl1_22
rlabel metal1 s 14094 0 14130 395 4 br1_22
rlabel metal1 s 14862 0 14898 395 4 bl0_23
rlabel metal1 s 14790 0 14826 395 4 br0_23
rlabel metal1 s 14646 0 14682 395 4 bl1_23
rlabel metal1 s 14574 0 14610 395 4 br1_23
rlabel metal1 s 15054 0 15090 395 4 bl0_24
rlabel metal1 s 15126 0 15162 395 4 br0_24
rlabel metal1 s 15270 0 15306 395 4 bl1_24
rlabel metal1 s 15342 0 15378 395 4 br1_24
rlabel metal1 s 16110 0 16146 395 4 bl0_25
rlabel metal1 s 16038 0 16074 395 4 br0_25
rlabel metal1 s 15894 0 15930 395 4 bl1_25
rlabel metal1 s 15822 0 15858 395 4 br1_25
rlabel metal1 s 16302 0 16338 395 4 bl0_26
rlabel metal1 s 16374 0 16410 395 4 br0_26
rlabel metal1 s 16518 0 16554 395 4 bl1_26
rlabel metal1 s 16590 0 16626 395 4 br1_26
rlabel metal1 s 17358 0 17394 395 4 bl0_27
rlabel metal1 s 17286 0 17322 395 4 br0_27
rlabel metal1 s 17142 0 17178 395 4 bl1_27
rlabel metal1 s 17070 0 17106 395 4 br1_27
rlabel metal1 s 17550 0 17586 395 4 bl0_28
rlabel metal1 s 17622 0 17658 395 4 br0_28
rlabel metal1 s 17766 0 17802 395 4 bl1_28
rlabel metal1 s 17838 0 17874 395 4 br1_28
rlabel metal1 s 18606 0 18642 395 4 bl0_29
rlabel metal1 s 18534 0 18570 395 4 br0_29
rlabel metal1 s 18390 0 18426 395 4 bl1_29
rlabel metal1 s 18318 0 18354 395 4 br1_29
rlabel metal1 s 18798 0 18834 395 4 bl0_30
rlabel metal1 s 18870 0 18906 395 4 br0_30
rlabel metal1 s 19014 0 19050 395 4 bl1_30
rlabel metal1 s 19086 0 19122 395 4 br1_30
rlabel metal1 s 19854 0 19890 395 4 bl0_31
rlabel metal1 s 19782 0 19818 395 4 br0_31
rlabel metal1 s 19638 0 19674 395 4 bl1_31
rlabel metal1 s 19566 0 19602 395 4 br1_31
rlabel metal1 s 20046 0 20082 395 4 bl0_32
rlabel metal1 s 20118 0 20154 395 4 br0_32
rlabel metal1 s 20262 0 20298 395 4 bl1_32
rlabel metal1 s 20334 0 20370 395 4 br1_32
rlabel metal1 s 21102 0 21138 395 4 bl0_33
rlabel metal1 s 21030 0 21066 395 4 br0_33
rlabel metal1 s 20886 0 20922 395 4 bl1_33
rlabel metal1 s 20814 0 20850 395 4 br1_33
rlabel metal1 s 21294 0 21330 395 4 bl0_34
rlabel metal1 s 21366 0 21402 395 4 br0_34
rlabel metal1 s 21510 0 21546 395 4 bl1_34
rlabel metal1 s 21582 0 21618 395 4 br1_34
rlabel metal1 s 22350 0 22386 395 4 bl0_35
rlabel metal1 s 22278 0 22314 395 4 br0_35
rlabel metal1 s 22134 0 22170 395 4 bl1_35
rlabel metal1 s 22062 0 22098 395 4 br1_35
rlabel metal1 s 22542 0 22578 395 4 bl0_36
rlabel metal1 s 22614 0 22650 395 4 br0_36
rlabel metal1 s 22758 0 22794 395 4 bl1_36
rlabel metal1 s 22830 0 22866 395 4 br1_36
rlabel metal1 s 23598 0 23634 395 4 bl0_37
rlabel metal1 s 23526 0 23562 395 4 br0_37
rlabel metal1 s 23382 0 23418 395 4 bl1_37
rlabel metal1 s 23310 0 23346 395 4 br1_37
rlabel metal1 s 23790 0 23826 395 4 bl0_38
rlabel metal1 s 23862 0 23898 395 4 br0_38
rlabel metal1 s 24006 0 24042 395 4 bl1_38
rlabel metal1 s 24078 0 24114 395 4 br1_38
rlabel metal1 s 24846 0 24882 395 4 bl0_39
rlabel metal1 s 24774 0 24810 395 4 br0_39
rlabel metal1 s 24630 0 24666 395 4 bl1_39
rlabel metal1 s 24558 0 24594 395 4 br1_39
rlabel metal1 s 25038 0 25074 395 4 bl0_40
rlabel metal1 s 25110 0 25146 395 4 br0_40
rlabel metal1 s 25254 0 25290 395 4 bl1_40
rlabel metal1 s 25326 0 25362 395 4 br1_40
rlabel metal1 s 26094 0 26130 395 4 bl0_41
rlabel metal1 s 26022 0 26058 395 4 br0_41
rlabel metal1 s 25878 0 25914 395 4 bl1_41
rlabel metal1 s 25806 0 25842 395 4 br1_41
rlabel metal1 s 26286 0 26322 395 4 bl0_42
rlabel metal1 s 26358 0 26394 395 4 br0_42
rlabel metal1 s 26502 0 26538 395 4 bl1_42
rlabel metal1 s 26574 0 26610 395 4 br1_42
rlabel metal1 s 27342 0 27378 395 4 bl0_43
rlabel metal1 s 27270 0 27306 395 4 br0_43
rlabel metal1 s 27126 0 27162 395 4 bl1_43
rlabel metal1 s 27054 0 27090 395 4 br1_43
rlabel metal1 s 27534 0 27570 395 4 bl0_44
rlabel metal1 s 27606 0 27642 395 4 br0_44
rlabel metal1 s 27750 0 27786 395 4 bl1_44
rlabel metal1 s 27822 0 27858 395 4 br1_44
rlabel metal1 s 28590 0 28626 395 4 bl0_45
rlabel metal1 s 28518 0 28554 395 4 br0_45
rlabel metal1 s 28374 0 28410 395 4 bl1_45
rlabel metal1 s 28302 0 28338 395 4 br1_45
rlabel metal1 s 28782 0 28818 395 4 bl0_46
rlabel metal1 s 28854 0 28890 395 4 br0_46
rlabel metal1 s 28998 0 29034 395 4 bl1_46
rlabel metal1 s 29070 0 29106 395 4 br1_46
rlabel metal1 s 29838 0 29874 395 4 bl0_47
rlabel metal1 s 29766 0 29802 395 4 br0_47
rlabel metal1 s 29622 0 29658 395 4 bl1_47
rlabel metal1 s 29550 0 29586 395 4 br1_47
rlabel metal1 s 30030 0 30066 395 4 bl0_48
rlabel metal1 s 30102 0 30138 395 4 br0_48
rlabel metal1 s 30246 0 30282 395 4 bl1_48
rlabel metal1 s 30318 0 30354 395 4 br1_48
rlabel metal1 s 31086 0 31122 395 4 bl0_49
rlabel metal1 s 31014 0 31050 395 4 br0_49
rlabel metal1 s 30870 0 30906 395 4 bl1_49
rlabel metal1 s 30798 0 30834 395 4 br1_49
rlabel metal1 s 31278 0 31314 395 4 bl0_50
rlabel metal1 s 31350 0 31386 395 4 br0_50
rlabel metal1 s 31494 0 31530 395 4 bl1_50
rlabel metal1 s 31566 0 31602 395 4 br1_50
rlabel metal1 s 32334 0 32370 395 4 bl0_51
rlabel metal1 s 32262 0 32298 395 4 br0_51
rlabel metal1 s 32118 0 32154 395 4 bl1_51
rlabel metal1 s 32046 0 32082 395 4 br1_51
rlabel metal1 s 32526 0 32562 395 4 bl0_52
rlabel metal1 s 32598 0 32634 395 4 br0_52
rlabel metal1 s 32742 0 32778 395 4 bl1_52
rlabel metal1 s 32814 0 32850 395 4 br1_52
rlabel metal1 s 33582 0 33618 395 4 bl0_53
rlabel metal1 s 33510 0 33546 395 4 br0_53
rlabel metal1 s 33366 0 33402 395 4 bl1_53
rlabel metal1 s 33294 0 33330 395 4 br1_53
rlabel metal1 s 33774 0 33810 395 4 bl0_54
rlabel metal1 s 33846 0 33882 395 4 br0_54
rlabel metal1 s 33990 0 34026 395 4 bl1_54
rlabel metal1 s 34062 0 34098 395 4 br1_54
rlabel metal1 s 34830 0 34866 395 4 bl0_55
rlabel metal1 s 34758 0 34794 395 4 br0_55
rlabel metal1 s 34614 0 34650 395 4 bl1_55
rlabel metal1 s 34542 0 34578 395 4 br1_55
rlabel metal1 s 35022 0 35058 395 4 bl0_56
rlabel metal1 s 35094 0 35130 395 4 br0_56
rlabel metal1 s 35238 0 35274 395 4 bl1_56
rlabel metal1 s 35310 0 35346 395 4 br1_56
rlabel metal1 s 36078 0 36114 395 4 bl0_57
rlabel metal1 s 36006 0 36042 395 4 br0_57
rlabel metal1 s 35862 0 35898 395 4 bl1_57
rlabel metal1 s 35790 0 35826 395 4 br1_57
rlabel metal1 s 36270 0 36306 395 4 bl0_58
rlabel metal1 s 36342 0 36378 395 4 br0_58
rlabel metal1 s 36486 0 36522 395 4 bl1_58
rlabel metal1 s 36558 0 36594 395 4 br1_58
rlabel metal1 s 37326 0 37362 395 4 bl0_59
rlabel metal1 s 37254 0 37290 395 4 br0_59
rlabel metal1 s 37110 0 37146 395 4 bl1_59
rlabel metal1 s 37038 0 37074 395 4 br1_59
rlabel metal1 s 37518 0 37554 395 4 bl0_60
rlabel metal1 s 37590 0 37626 395 4 br0_60
rlabel metal1 s 37734 0 37770 395 4 bl1_60
rlabel metal1 s 37806 0 37842 395 4 br1_60
rlabel metal1 s 38574 0 38610 395 4 bl0_61
rlabel metal1 s 38502 0 38538 395 4 br0_61
rlabel metal1 s 38358 0 38394 395 4 bl1_61
rlabel metal1 s 38286 0 38322 395 4 br1_61
rlabel metal1 s 38766 0 38802 395 4 bl0_62
rlabel metal1 s 38838 0 38874 395 4 br0_62
rlabel metal1 s 38982 0 39018 395 4 bl1_62
rlabel metal1 s 39054 0 39090 395 4 br1_62
rlabel metal1 s 39822 0 39858 395 4 bl0_63
rlabel metal1 s 39750 0 39786 395 4 br0_63
rlabel metal1 s 39606 0 39642 395 4 bl1_63
rlabel metal1 s 39534 0 39570 395 4 br1_63
rlabel metal1 s 40014 0 40050 395 4 bl0_64
rlabel metal1 s 40086 0 40122 395 4 br0_64
rlabel metal1 s 40230 0 40266 395 4 bl1_64
rlabel metal1 s 40302 0 40338 395 4 br1_64
rlabel metal1 s 41070 0 41106 395 4 bl0_65
rlabel metal1 s 40998 0 41034 395 4 br0_65
rlabel metal1 s 40854 0 40890 395 4 bl1_65
rlabel metal1 s 40782 0 40818 395 4 br1_65
rlabel metal1 s 41262 0 41298 395 4 bl0_66
rlabel metal1 s 41334 0 41370 395 4 br0_66
rlabel metal1 s 41478 0 41514 395 4 bl1_66
rlabel metal1 s 41550 0 41586 395 4 br1_66
rlabel metal1 s 42318 0 42354 395 4 bl0_67
rlabel metal1 s 42246 0 42282 395 4 br0_67
rlabel metal1 s 42102 0 42138 395 4 bl1_67
rlabel metal1 s 42030 0 42066 395 4 br1_67
rlabel metal1 s 42510 0 42546 395 4 bl0_68
rlabel metal1 s 42582 0 42618 395 4 br0_68
rlabel metal1 s 42726 0 42762 395 4 bl1_68
rlabel metal1 s 42798 0 42834 395 4 br1_68
rlabel metal1 s 43566 0 43602 395 4 bl0_69
rlabel metal1 s 43494 0 43530 395 4 br0_69
rlabel metal1 s 43350 0 43386 395 4 bl1_69
rlabel metal1 s 43278 0 43314 395 4 br1_69
rlabel metal1 s 43758 0 43794 395 4 bl0_70
rlabel metal1 s 43830 0 43866 395 4 br0_70
rlabel metal1 s 43974 0 44010 395 4 bl1_70
rlabel metal1 s 44046 0 44082 395 4 br1_70
rlabel metal1 s 44814 0 44850 395 4 bl0_71
rlabel metal1 s 44742 0 44778 395 4 br0_71
rlabel metal1 s 44598 0 44634 395 4 bl1_71
rlabel metal1 s 44526 0 44562 395 4 br1_71
rlabel metal1 s 45006 0 45042 395 4 bl0_72
rlabel metal1 s 45078 0 45114 395 4 br0_72
rlabel metal1 s 45222 0 45258 395 4 bl1_72
rlabel metal1 s 45294 0 45330 395 4 br1_72
rlabel metal1 s 46062 0 46098 395 4 bl0_73
rlabel metal1 s 45990 0 46026 395 4 br0_73
rlabel metal1 s 45846 0 45882 395 4 bl1_73
rlabel metal1 s 45774 0 45810 395 4 br1_73
rlabel metal1 s 46254 0 46290 395 4 bl0_74
rlabel metal1 s 46326 0 46362 395 4 br0_74
rlabel metal1 s 46470 0 46506 395 4 bl1_74
rlabel metal1 s 46542 0 46578 395 4 br1_74
rlabel metal1 s 47310 0 47346 395 4 bl0_75
rlabel metal1 s 47238 0 47274 395 4 br0_75
rlabel metal1 s 47094 0 47130 395 4 bl1_75
rlabel metal1 s 47022 0 47058 395 4 br1_75
rlabel metal1 s 47502 0 47538 395 4 bl0_76
rlabel metal1 s 47574 0 47610 395 4 br0_76
rlabel metal1 s 47718 0 47754 395 4 bl1_76
rlabel metal1 s 47790 0 47826 395 4 br1_76
rlabel metal1 s 48558 0 48594 395 4 bl0_77
rlabel metal1 s 48486 0 48522 395 4 br0_77
rlabel metal1 s 48342 0 48378 395 4 bl1_77
rlabel metal1 s 48270 0 48306 395 4 br1_77
rlabel metal1 s 48750 0 48786 395 4 bl0_78
rlabel metal1 s 48822 0 48858 395 4 br0_78
rlabel metal1 s 48966 0 49002 395 4 bl1_78
rlabel metal1 s 49038 0 49074 395 4 br1_78
rlabel metal1 s 49806 0 49842 395 4 bl0_79
rlabel metal1 s 49734 0 49770 395 4 br0_79
rlabel metal1 s 49590 0 49626 395 4 bl1_79
rlabel metal1 s 49518 0 49554 395 4 br1_79
rlabel metal1 s 49998 0 50034 395 4 bl0_80
rlabel metal1 s 50070 0 50106 395 4 br0_80
rlabel metal1 s 50214 0 50250 395 4 bl1_80
rlabel metal1 s 50286 0 50322 395 4 br1_80
rlabel metal1 s 51054 0 51090 395 4 bl0_81
rlabel metal1 s 50982 0 51018 395 4 br0_81
rlabel metal1 s 50838 0 50874 395 4 bl1_81
rlabel metal1 s 50766 0 50802 395 4 br1_81
rlabel metal1 s 51246 0 51282 395 4 bl0_82
rlabel metal1 s 51318 0 51354 395 4 br0_82
rlabel metal1 s 51462 0 51498 395 4 bl1_82
rlabel metal1 s 51534 0 51570 395 4 br1_82
rlabel metal1 s 52302 0 52338 395 4 bl0_83
rlabel metal1 s 52230 0 52266 395 4 br0_83
rlabel metal1 s 52086 0 52122 395 4 bl1_83
rlabel metal1 s 52014 0 52050 395 4 br1_83
rlabel metal1 s 52494 0 52530 395 4 bl0_84
rlabel metal1 s 52566 0 52602 395 4 br0_84
rlabel metal1 s 52710 0 52746 395 4 bl1_84
rlabel metal1 s 52782 0 52818 395 4 br1_84
rlabel metal1 s 53550 0 53586 395 4 bl0_85
rlabel metal1 s 53478 0 53514 395 4 br0_85
rlabel metal1 s 53334 0 53370 395 4 bl1_85
rlabel metal1 s 53262 0 53298 395 4 br1_85
rlabel metal1 s 53742 0 53778 395 4 bl0_86
rlabel metal1 s 53814 0 53850 395 4 br0_86
rlabel metal1 s 53958 0 53994 395 4 bl1_86
rlabel metal1 s 54030 0 54066 395 4 br1_86
rlabel metal1 s 54798 0 54834 395 4 bl0_87
rlabel metal1 s 54726 0 54762 395 4 br0_87
rlabel metal1 s 54582 0 54618 395 4 bl1_87
rlabel metal1 s 54510 0 54546 395 4 br1_87
rlabel metal1 s 54990 0 55026 395 4 bl0_88
rlabel metal1 s 55062 0 55098 395 4 br0_88
rlabel metal1 s 55206 0 55242 395 4 bl1_88
rlabel metal1 s 55278 0 55314 395 4 br1_88
rlabel metal1 s 56046 0 56082 395 4 bl0_89
rlabel metal1 s 55974 0 56010 395 4 br0_89
rlabel metal1 s 55830 0 55866 395 4 bl1_89
rlabel metal1 s 55758 0 55794 395 4 br1_89
rlabel metal1 s 56238 0 56274 395 4 bl0_90
rlabel metal1 s 56310 0 56346 395 4 br0_90
rlabel metal1 s 56454 0 56490 395 4 bl1_90
rlabel metal1 s 56526 0 56562 395 4 br1_90
rlabel metal1 s 57294 0 57330 395 4 bl0_91
rlabel metal1 s 57222 0 57258 395 4 br0_91
rlabel metal1 s 57078 0 57114 395 4 bl1_91
rlabel metal1 s 57006 0 57042 395 4 br1_91
rlabel metal1 s 57486 0 57522 395 4 bl0_92
rlabel metal1 s 57558 0 57594 395 4 br0_92
rlabel metal1 s 57702 0 57738 395 4 bl1_92
rlabel metal1 s 57774 0 57810 395 4 br1_92
rlabel metal1 s 58542 0 58578 395 4 bl0_93
rlabel metal1 s 58470 0 58506 395 4 br0_93
rlabel metal1 s 58326 0 58362 395 4 bl1_93
rlabel metal1 s 58254 0 58290 395 4 br1_93
rlabel metal1 s 58734 0 58770 395 4 bl0_94
rlabel metal1 s 58806 0 58842 395 4 br0_94
rlabel metal1 s 58950 0 58986 395 4 bl1_94
rlabel metal1 s 59022 0 59058 395 4 br1_94
rlabel metal1 s 59790 0 59826 395 4 bl0_95
rlabel metal1 s 59718 0 59754 395 4 br0_95
rlabel metal1 s 59574 0 59610 395 4 bl1_95
rlabel metal1 s 59502 0 59538 395 4 br1_95
rlabel metal1 s 59982 0 60018 395 4 bl0_96
rlabel metal1 s 60054 0 60090 395 4 br0_96
rlabel metal1 s 60198 0 60234 395 4 bl1_96
rlabel metal1 s 60270 0 60306 395 4 br1_96
rlabel metal1 s 61038 0 61074 395 4 bl0_97
rlabel metal1 s 60966 0 61002 395 4 br0_97
rlabel metal1 s 60822 0 60858 395 4 bl1_97
rlabel metal1 s 60750 0 60786 395 4 br1_97
rlabel metal1 s 61230 0 61266 395 4 bl0_98
rlabel metal1 s 61302 0 61338 395 4 br0_98
rlabel metal1 s 61446 0 61482 395 4 bl1_98
rlabel metal1 s 61518 0 61554 395 4 br1_98
rlabel metal1 s 62286 0 62322 395 4 bl0_99
rlabel metal1 s 62214 0 62250 395 4 br0_99
rlabel metal1 s 62070 0 62106 395 4 bl1_99
rlabel metal1 s 61998 0 62034 395 4 br1_99
rlabel metal1 s 62478 0 62514 395 4 bl0_100
rlabel metal1 s 62550 0 62586 395 4 br0_100
rlabel metal1 s 62694 0 62730 395 4 bl1_100
rlabel metal1 s 62766 0 62802 395 4 br1_100
rlabel metal1 s 63534 0 63570 395 4 bl0_101
rlabel metal1 s 63462 0 63498 395 4 br0_101
rlabel metal1 s 63318 0 63354 395 4 bl1_101
rlabel metal1 s 63246 0 63282 395 4 br1_101
rlabel metal1 s 63726 0 63762 395 4 bl0_102
rlabel metal1 s 63798 0 63834 395 4 br0_102
rlabel metal1 s 63942 0 63978 395 4 bl1_102
rlabel metal1 s 64014 0 64050 395 4 br1_102
rlabel metal1 s 64782 0 64818 395 4 bl0_103
rlabel metal1 s 64710 0 64746 395 4 br0_103
rlabel metal1 s 64566 0 64602 395 4 bl1_103
rlabel metal1 s 64494 0 64530 395 4 br1_103
rlabel metal1 s 64974 0 65010 395 4 bl0_104
rlabel metal1 s 65046 0 65082 395 4 br0_104
rlabel metal1 s 65190 0 65226 395 4 bl1_104
rlabel metal1 s 65262 0 65298 395 4 br1_104
rlabel metal1 s 66030 0 66066 395 4 bl0_105
rlabel metal1 s 65958 0 65994 395 4 br0_105
rlabel metal1 s 65814 0 65850 395 4 bl1_105
rlabel metal1 s 65742 0 65778 395 4 br1_105
rlabel metal1 s 66222 0 66258 395 4 bl0_106
rlabel metal1 s 66294 0 66330 395 4 br0_106
rlabel metal1 s 66438 0 66474 395 4 bl1_106
rlabel metal1 s 66510 0 66546 395 4 br1_106
rlabel metal1 s 67278 0 67314 395 4 bl0_107
rlabel metal1 s 67206 0 67242 395 4 br0_107
rlabel metal1 s 67062 0 67098 395 4 bl1_107
rlabel metal1 s 66990 0 67026 395 4 br1_107
rlabel metal1 s 67470 0 67506 395 4 bl0_108
rlabel metal1 s 67542 0 67578 395 4 br0_108
rlabel metal1 s 67686 0 67722 395 4 bl1_108
rlabel metal1 s 67758 0 67794 395 4 br1_108
rlabel metal1 s 68526 0 68562 395 4 bl0_109
rlabel metal1 s 68454 0 68490 395 4 br0_109
rlabel metal1 s 68310 0 68346 395 4 bl1_109
rlabel metal1 s 68238 0 68274 395 4 br1_109
rlabel metal1 s 68718 0 68754 395 4 bl0_110
rlabel metal1 s 68790 0 68826 395 4 br0_110
rlabel metal1 s 68934 0 68970 395 4 bl1_110
rlabel metal1 s 69006 0 69042 395 4 br1_110
rlabel metal1 s 69774 0 69810 395 4 bl0_111
rlabel metal1 s 69702 0 69738 395 4 br0_111
rlabel metal1 s 69558 0 69594 395 4 bl1_111
rlabel metal1 s 69486 0 69522 395 4 br1_111
rlabel metal1 s 69966 0 70002 395 4 bl0_112
rlabel metal1 s 70038 0 70074 395 4 br0_112
rlabel metal1 s 70182 0 70218 395 4 bl1_112
rlabel metal1 s 70254 0 70290 395 4 br1_112
rlabel metal1 s 71022 0 71058 395 4 bl0_113
rlabel metal1 s 70950 0 70986 395 4 br0_113
rlabel metal1 s 70806 0 70842 395 4 bl1_113
rlabel metal1 s 70734 0 70770 395 4 br1_113
rlabel metal1 s 71214 0 71250 395 4 bl0_114
rlabel metal1 s 71286 0 71322 395 4 br0_114
rlabel metal1 s 71430 0 71466 395 4 bl1_114
rlabel metal1 s 71502 0 71538 395 4 br1_114
rlabel metal1 s 72270 0 72306 395 4 bl0_115
rlabel metal1 s 72198 0 72234 395 4 br0_115
rlabel metal1 s 72054 0 72090 395 4 bl1_115
rlabel metal1 s 71982 0 72018 395 4 br1_115
rlabel metal1 s 72462 0 72498 395 4 bl0_116
rlabel metal1 s 72534 0 72570 395 4 br0_116
rlabel metal1 s 72678 0 72714 395 4 bl1_116
rlabel metal1 s 72750 0 72786 395 4 br1_116
rlabel metal1 s 73518 0 73554 395 4 bl0_117
rlabel metal1 s 73446 0 73482 395 4 br0_117
rlabel metal1 s 73302 0 73338 395 4 bl1_117
rlabel metal1 s 73230 0 73266 395 4 br1_117
rlabel metal1 s 73710 0 73746 395 4 bl0_118
rlabel metal1 s 73782 0 73818 395 4 br0_118
rlabel metal1 s 73926 0 73962 395 4 bl1_118
rlabel metal1 s 73998 0 74034 395 4 br1_118
rlabel metal1 s 74766 0 74802 395 4 bl0_119
rlabel metal1 s 74694 0 74730 395 4 br0_119
rlabel metal1 s 74550 0 74586 395 4 bl1_119
rlabel metal1 s 74478 0 74514 395 4 br1_119
rlabel metal1 s 74958 0 74994 395 4 bl0_120
rlabel metal1 s 75030 0 75066 395 4 br0_120
rlabel metal1 s 75174 0 75210 395 4 bl1_120
rlabel metal1 s 75246 0 75282 395 4 br1_120
rlabel metal1 s 76014 0 76050 395 4 bl0_121
rlabel metal1 s 75942 0 75978 395 4 br0_121
rlabel metal1 s 75798 0 75834 395 4 bl1_121
rlabel metal1 s 75726 0 75762 395 4 br1_121
rlabel metal1 s 76206 0 76242 395 4 bl0_122
rlabel metal1 s 76278 0 76314 395 4 br0_122
rlabel metal1 s 76422 0 76458 395 4 bl1_122
rlabel metal1 s 76494 0 76530 395 4 br1_122
rlabel metal1 s 77262 0 77298 395 4 bl0_123
rlabel metal1 s 77190 0 77226 395 4 br0_123
rlabel metal1 s 77046 0 77082 395 4 bl1_123
rlabel metal1 s 76974 0 77010 395 4 br1_123
rlabel metal1 s 77454 0 77490 395 4 bl0_124
rlabel metal1 s 77526 0 77562 395 4 br0_124
rlabel metal1 s 77670 0 77706 395 4 bl1_124
rlabel metal1 s 77742 0 77778 395 4 br1_124
rlabel metal1 s 78510 0 78546 395 4 bl0_125
rlabel metal1 s 78438 0 78474 395 4 br0_125
rlabel metal1 s 78294 0 78330 395 4 bl1_125
rlabel metal1 s 78222 0 78258 395 4 br1_125
rlabel metal1 s 78702 0 78738 395 4 bl0_126
rlabel metal1 s 78774 0 78810 395 4 br0_126
rlabel metal1 s 78918 0 78954 395 4 bl1_126
rlabel metal1 s 78990 0 79026 395 4 br1_126
rlabel metal1 s 79758 0 79794 395 4 bl0_127
rlabel metal1 s 79686 0 79722 395 4 br0_127
rlabel metal1 s 79542 0 79578 395 4 bl1_127
rlabel metal1 s 79470 0 79506 395 4 br1_127
<< properties >>
string FIXED_BBOX 0 0 79872 474
string GDS_END 1959538
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 1827342
<< end >>
