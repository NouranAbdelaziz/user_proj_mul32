magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal3 >>
rect 106 11282 4879 11346
rect 10078 11282 14858 11346
rect 10078 10330 14858 10564
rect 106 9548 4879 9612
rect 10078 9548 14858 9612
rect 194 7348 4879 8036
rect 10078 7348 14858 8036
<< obsm3 >>
rect 99 10330 4879 10564
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 4874 11347
rect 10083 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 4874 10565
rect 14746 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 4874 9613
rect 10083 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 4874 8037
rect 10083 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< obsm4 >>
rect 334 35077 14666 40000
rect 193 19080 14807 35077
rect 334 13927 14666 19080
rect 193 13787 14807 13927
rect 334 12737 14666 13787
rect 193 12617 14807 12737
rect 334 11567 14666 12617
rect 193 11427 14807 11567
rect 4954 11301 10003 11427
rect 4954 10349 14666 10545
rect 4954 9467 10003 9593
rect 193 9327 14807 9467
rect 334 8237 14666 9327
rect 193 8117 14807 8237
rect 4954 7267 10003 8117
rect 193 7147 14807 7267
rect 334 6297 14666 7147
rect 193 6177 14807 6297
rect 334 5087 14666 6177
rect 193 4967 14807 5087
rect 334 3877 14666 4967
rect 193 3757 14807 3877
rect 273 2907 14727 3757
rect 193 2787 14807 2907
rect 334 1697 14666 2787
rect 193 1577 14807 1697
rect 334 407 14666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 574 34837 14426 40000
rect 0 19317 15000 34837
rect 574 7368 14426 19317
rect 0 7367 15000 7368
rect 574 3657 14426 7367
rect 513 3007 14487 3657
rect 574 427 14426 3007
<< labels >>
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 10625 254 11221 6 AMUXBUS_A
port 2 nsew signal bidirectional
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 2 nsew signal bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 3 nsew signal bidirectional
rlabel metal4 s 0 9673 254 10269 6 AMUXBUS_B
port 4 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 4 nsew signal bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 5 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 6 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 12 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 12 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 12 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 12 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 13 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 14 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 15 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 16 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 16 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 16 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 16 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 17 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 18 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 19 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 20 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 21 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 22 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 23 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 24 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 24 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 24 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 25 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 26 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 27 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 28 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 28 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 28 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 28 nsew power bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 29 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 31 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 32 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 33 nsew ground bidirectional
rlabel metal4 s 0 9547 254 9613 6 VSSA
port 34 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 35 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 6 VSSA
port 36 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 37 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 38 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 106 9548 4879 9612 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 106 11282 4879 11346 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 194 7348 4879 8036 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10078 7348 14858 8036 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10078 9548 14858 9612 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10078 10330 14858 10564 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10078 11282 14858 11346 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 0 7347 4874 8037 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 0 9547 4874 9613 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 0 10329 4874 10565 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 0 11281 4874 11347 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 10083 7347 15000 8037 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 10083 9547 15000 9613 6 VSSA
port 40 nsew ground bidirectional
rlabel metal4 s 10083 11281 15000 11347 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 11294 14840 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 10511 14840 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 10427 14840 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 10343 14840 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 9560 14840 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 7980 14840 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 7892 14840 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 7804 14840 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 7716 14840 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 7628 14840 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 7540 14840 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 7452 14840 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14800 7364 14840 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 10511 14759 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 10427 14759 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 10343 14759 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 7980 14759 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 7892 14759 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 7804 14759 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 7716 14759 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 7628 14759 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 7540 14759 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 7452 14759 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14719 7364 14759 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14718 11294 14758 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14718 9560 14758 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 10511 14678 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 10427 14678 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 10343 14678 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 7980 14678 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 7892 14678 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 7804 14678 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 7716 14678 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 7628 14678 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 7540 14678 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 7452 14678 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14638 7364 14678 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14636 11294 14676 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14636 9560 14676 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 10511 14597 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 10427 14597 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 10343 14597 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 7980 14597 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 7892 14597 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 7804 14597 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 7716 14597 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 7628 14597 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 7540 14597 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 7452 14597 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14557 7364 14597 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14554 11294 14594 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14554 9560 14594 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 10511 14516 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 10427 14516 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 10343 14516 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 7980 14516 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 7892 14516 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 7804 14516 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 7716 14516 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 7628 14516 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 7540 14516 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 7452 14516 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14476 7364 14516 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14472 11294 14512 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14472 9560 14512 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 10511 14435 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 10427 14435 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 10343 14435 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 7980 14435 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 7892 14435 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 7804 14435 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 7716 14435 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 7628 14435 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 7540 14435 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 7452 14435 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14395 7364 14435 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14390 11294 14430 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14390 9560 14430 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 10511 14354 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 10427 14354 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 10343 14354 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 7980 14354 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 7892 14354 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 7804 14354 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 7716 14354 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 7628 14354 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 7540 14354 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 7452 14354 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14314 7364 14354 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14308 11294 14348 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14308 9560 14348 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 10511 14273 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 10427 14273 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 10343 14273 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 7980 14273 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 7892 14273 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 7804 14273 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 7716 14273 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 7628 14273 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 7540 14273 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 7452 14273 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14233 7364 14273 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14227 11294 14267 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14227 9560 14267 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 10511 14192 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 10427 14192 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 10343 14192 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 7980 14192 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 7892 14192 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 7804 14192 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 7716 14192 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 7628 14192 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 7540 14192 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 7452 14192 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14152 7364 14192 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14146 11294 14186 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14146 9560 14186 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 10511 14111 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 10427 14111 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 10343 14111 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 7980 14111 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 7892 14111 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 7804 14111 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 7716 14111 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 7628 14111 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 7540 14111 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 7452 14111 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14071 7364 14111 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14065 11294 14105 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 14065 9560 14105 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 10511 14030 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 10427 14030 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 10343 14030 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 7980 14030 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 7892 14030 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 7804 14030 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 7716 14030 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 7628 14030 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 7540 14030 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 7452 14030 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13990 7364 14030 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13984 11294 14024 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13984 9560 14024 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 10511 13949 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 10427 13949 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 10343 13949 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 7980 13949 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 7892 13949 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 7804 13949 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 7716 13949 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 7628 13949 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 7540 13949 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 7452 13949 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13909 7364 13949 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13903 11294 13943 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13903 9560 13943 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 10511 13868 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 10427 13868 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 10343 13868 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 7980 13868 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 7892 13868 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 7804 13868 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 7716 13868 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 7628 13868 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 7540 13868 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 7452 13868 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13828 7364 13868 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13822 11294 13862 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13822 9560 13862 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 10511 13787 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 10427 13787 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 10343 13787 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 7980 13787 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 7892 13787 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 7804 13787 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 7716 13787 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 7628 13787 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 7540 13787 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 7452 13787 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13747 7364 13787 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13741 11294 13781 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13741 9560 13781 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 10511 13706 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 10427 13706 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 10343 13706 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 7980 13706 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 7892 13706 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 7804 13706 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 7716 13706 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 7628 13706 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 7540 13706 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 7452 13706 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13666 7364 13706 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13660 11294 13700 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13660 9560 13700 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 10511 13625 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 10427 13625 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 10343 13625 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 7980 13625 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 7892 13625 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 7804 13625 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 7716 13625 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 7628 13625 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 7540 13625 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 7452 13625 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13585 7364 13625 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13579 11294 13619 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13579 9560 13619 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 10511 13544 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 10427 13544 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 10343 13544 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 7980 13544 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 7892 13544 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 7804 13544 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 7716 13544 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 7628 13544 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 7540 13544 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 7452 13544 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13504 7364 13544 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13498 11294 13538 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13498 9560 13538 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 10511 13463 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 10427 13463 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 10343 13463 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 7980 13463 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 7892 13463 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 7804 13463 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 7716 13463 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 7628 13463 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 7540 13463 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 7452 13463 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13423 7364 13463 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13417 11294 13457 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13417 9560 13457 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 10511 13382 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 10427 13382 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 10343 13382 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 7980 13382 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 7892 13382 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 7804 13382 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 7716 13382 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 7628 13382 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 7540 13382 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 7452 13382 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13342 7364 13382 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13336 11294 13376 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13336 9560 13376 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 10511 13301 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 10427 13301 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 10343 13301 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 7980 13301 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 7892 13301 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 7804 13301 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 7716 13301 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 7628 13301 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 7540 13301 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 7452 13301 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13261 7364 13301 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13255 11294 13295 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13255 9560 13295 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 10511 13220 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 10427 13220 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 10343 13220 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 7980 13220 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 7892 13220 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 7804 13220 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 7716 13220 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 7628 13220 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 7540 13220 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 7452 13220 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13180 7364 13220 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13174 11294 13214 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13174 9560 13214 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 10511 13139 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 10427 13139 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 10343 13139 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 7980 13139 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 7892 13139 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 7804 13139 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 7716 13139 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 7628 13139 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 7540 13139 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 7452 13139 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13099 7364 13139 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13093 11294 13133 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13093 9560 13133 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 10511 13058 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 10427 13058 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 10343 13058 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 7980 13058 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 7892 13058 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 7804 13058 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 7716 13058 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 7628 13058 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 7540 13058 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 7452 13058 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13018 7364 13058 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13012 11294 13052 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 13012 9560 13052 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 10511 12977 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 10427 12977 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 10343 12977 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 7980 12977 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 7892 12977 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 7804 12977 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 7716 12977 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 7628 12977 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 7540 12977 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 7452 12977 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12937 7364 12977 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12931 11294 12971 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12931 9560 12971 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 10511 12896 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 10427 12896 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 10343 12896 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 7980 12896 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 7892 12896 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 7804 12896 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 7716 12896 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 7628 12896 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 7540 12896 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 7452 12896 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12856 7364 12896 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12850 11294 12890 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12850 9560 12890 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 10511 12815 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 10427 12815 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 10343 12815 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 7980 12815 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 7892 12815 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 7804 12815 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 7716 12815 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 7628 12815 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 7540 12815 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 7452 12815 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12775 7364 12815 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12769 11294 12809 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12769 9560 12809 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 10511 12734 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 10427 12734 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 10343 12734 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 7980 12734 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 7892 12734 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 7804 12734 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 7716 12734 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 7628 12734 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 7540 12734 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 7452 12734 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12694 7364 12734 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12688 11294 12728 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12688 9560 12728 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 10511 12653 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 10427 12653 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 10343 12653 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 7980 12653 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 7892 12653 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 7804 12653 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 7716 12653 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 7628 12653 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 7540 12653 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 7452 12653 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12613 7364 12653 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12607 11294 12647 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12607 9560 12647 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 10511 12572 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 10427 12572 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 10343 12572 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 7980 12572 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 7892 12572 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 7804 12572 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 7716 12572 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 7628 12572 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 7540 12572 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 7452 12572 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12532 7364 12572 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12526 11294 12566 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12526 9560 12566 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 10511 12491 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 10427 12491 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 10343 12491 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 7980 12491 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 7892 12491 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 7804 12491 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 7716 12491 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 7628 12491 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 7540 12491 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 7452 12491 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12451 7364 12491 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12445 11294 12485 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12445 9560 12485 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 10511 12410 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 10427 12410 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 10343 12410 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 7980 12410 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 7892 12410 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 7804 12410 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 7716 12410 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 7628 12410 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 7540 12410 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 7452 12410 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12370 7364 12410 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12364 11294 12404 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12364 9560 12404 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 10511 12329 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 10427 12329 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 10343 12329 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 7980 12329 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 7892 12329 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 7804 12329 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 7716 12329 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 7628 12329 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 7540 12329 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 7452 12329 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12289 7364 12329 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12283 11294 12323 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12283 9560 12323 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 10511 12248 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 10427 12248 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 10343 12248 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 7980 12248 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 7892 12248 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 7804 12248 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 7716 12248 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 7628 12248 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 7540 12248 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 7452 12248 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12208 7364 12248 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12202 11294 12242 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12202 9560 12242 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 10511 12167 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 10427 12167 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 10343 12167 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 7980 12167 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 7892 12167 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 7804 12167 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 7716 12167 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 7628 12167 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 7540 12167 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 7452 12167 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12127 7364 12167 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12121 11294 12161 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12121 9560 12161 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 10511 12086 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 10427 12086 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 10343 12086 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 7980 12086 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 7892 12086 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 7804 12086 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 7716 12086 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 7628 12086 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 7540 12086 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 7452 12086 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12046 7364 12086 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12040 11294 12080 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 12040 9560 12080 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 10511 12005 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 10427 12005 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 10343 12005 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 7980 12005 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 7892 12005 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 7804 12005 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 7716 12005 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 7628 12005 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 7540 12005 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 7452 12005 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11965 7364 12005 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11959 11294 11999 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11959 9560 11999 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 10511 11924 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 10427 11924 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 10343 11924 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 7980 11924 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 7892 11924 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 7804 11924 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 7716 11924 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 7628 11924 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 7540 11924 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 7452 11924 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11884 7364 11924 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11878 11294 11918 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11878 9560 11918 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 10511 11843 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 10427 11843 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 10343 11843 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 7980 11843 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 7892 11843 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 7804 11843 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 7716 11843 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 7628 11843 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 7540 11843 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 7452 11843 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11803 7364 11843 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11797 11294 11837 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11797 9560 11837 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 10511 11762 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 10427 11762 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 10343 11762 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 7980 11762 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 7892 11762 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 7804 11762 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 7716 11762 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 7628 11762 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 7540 11762 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 7452 11762 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11722 7364 11762 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11716 11294 11756 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11716 9560 11756 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 10511 11681 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 10427 11681 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 10343 11681 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 7980 11681 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 7892 11681 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 7804 11681 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 7716 11681 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 7628 11681 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 7540 11681 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 7452 11681 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11641 7364 11681 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11635 11294 11675 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11635 9560 11675 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 10511 11600 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 10427 11600 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 10343 11600 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 7980 11600 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 7892 11600 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 7804 11600 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 7716 11600 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 7628 11600 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 7540 11600 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 7452 11600 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11560 7364 11600 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11554 11294 11594 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11554 9560 11594 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 10511 11519 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 10427 11519 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 10343 11519 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 7980 11519 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 7892 11519 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 7804 11519 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 7716 11519 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 7628 11519 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 7540 11519 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 7452 11519 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11479 7364 11519 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11473 11294 11513 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11473 9560 11513 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 10511 11438 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 10427 11438 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 10343 11438 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 7980 11438 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 7892 11438 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 7804 11438 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 7716 11438 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 7628 11438 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 7540 11438 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 7452 11438 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11398 7364 11438 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11392 11294 11432 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11392 9560 11432 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 10511 11357 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 10427 11357 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 10343 11357 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 7980 11357 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 7892 11357 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 7804 11357 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 7716 11357 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 7628 11357 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 7540 11357 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 7452 11357 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11317 7364 11357 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11311 11294 11351 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11311 9560 11351 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 10511 11276 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 10427 11276 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 10343 11276 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 7980 11276 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 7892 11276 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 7804 11276 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 7716 11276 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 7628 11276 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 7540 11276 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 7452 11276 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11236 7364 11276 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11230 11294 11270 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11230 9560 11270 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 10511 11195 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 10427 11195 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 10343 11195 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 7980 11195 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 7892 11195 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 7804 11195 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 7716 11195 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 7628 11195 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 7540 11195 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 7452 11195 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11155 7364 11195 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11149 11294 11189 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11149 9560 11189 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 10511 11114 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 10427 11114 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 10343 11114 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 7980 11114 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 7892 11114 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 7804 11114 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 7716 11114 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 7628 11114 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 7540 11114 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 7452 11114 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11074 7364 11114 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11068 11294 11108 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 11068 9560 11108 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 10511 11033 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 10427 11033 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 10343 11033 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 7980 11033 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 7892 11033 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 7804 11033 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 7716 11033 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 7628 11033 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 7540 11033 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 7452 11033 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10993 7364 11033 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10987 11294 11027 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10987 9560 11027 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 10511 10952 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 10427 10952 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 10343 10952 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 7980 10952 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 7892 10952 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 7804 10952 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 7716 10952 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 7628 10952 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 7540 10952 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 7452 10952 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10912 7364 10952 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10906 11294 10946 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10906 9560 10946 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 10511 10871 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 10427 10871 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 10343 10871 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 7980 10871 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 7892 10871 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 7804 10871 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 7716 10871 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 7628 10871 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 7540 10871 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 7452 10871 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10831 7364 10871 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10825 11294 10865 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10825 9560 10865 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 10511 10790 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 10427 10790 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 10343 10790 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 7980 10790 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 7892 10790 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 7804 10790 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 7716 10790 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 7628 10790 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 7540 10790 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 7452 10790 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10750 7364 10790 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10744 11294 10784 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10744 9560 10784 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 10511 10709 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 10427 10709 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 10343 10709 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 7980 10709 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 7892 10709 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 7804 10709 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 7716 10709 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 7628 10709 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 7540 10709 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 7452 10709 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10669 7364 10709 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10663 11294 10703 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10663 9560 10703 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 10511 10628 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 10427 10628 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 10343 10628 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 7980 10628 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 7892 10628 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 7804 10628 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 7716 10628 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 7628 10628 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 7540 10628 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 7452 10628 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10588 7364 10628 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10582 11294 10622 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10582 9560 10622 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 10511 10546 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 10427 10546 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 10343 10546 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 7980 10546 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 7892 10546 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 7804 10546 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 7716 10546 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 7628 10546 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 7540 10546 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 7452 10546 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10506 7364 10546 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10501 11294 10541 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10501 9560 10541 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 10511 10464 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 10427 10464 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 10343 10464 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 7980 10464 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 7892 10464 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 7804 10464 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 7716 10464 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 7628 10464 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 7540 10464 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 7452 10464 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10424 7364 10464 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10420 11294 10460 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10420 9560 10460 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 10511 10382 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 10427 10382 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 10343 10382 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 7980 10382 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 7892 10382 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 7804 10382 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 7716 10382 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 7628 10382 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 7540 10382 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 7452 10382 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10342 7364 10382 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10339 11294 10379 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10339 9560 10379 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 10511 10300 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 10427 10300 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 10343 10300 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 7980 10300 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 7892 10300 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 7804 10300 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 7716 10300 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 7628 10300 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 7540 10300 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 7452 10300 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10260 7364 10300 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10258 11294 10298 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10258 9560 10298 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 10511 10218 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 10427 10218 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 10343 10218 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 7980 10218 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 7892 10218 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 7804 10218 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 7716 10218 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 7628 10218 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 7540 10218 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 7452 10218 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10178 7364 10218 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10177 11294 10217 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10177 9560 10217 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 11294 10136 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 10511 10136 10551 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 10427 10136 10467 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 10343 10136 10383 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 9560 10136 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 7980 10136 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 7892 10136 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 7804 10136 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 7716 10136 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 7628 10136 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 7540 10136 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 7452 10136 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 10096 7364 10136 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 11294 4861 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4809 10499 4873 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4809 10415 4873 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4809 10331 4873 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 9560 4861 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 7980 4861 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 7892 4861 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 7804 4861 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 7716 4861 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 7628 4861 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 7540 4861 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 7452 4861 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4821 7364 4861 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 11294 4781 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 9560 4781 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 7980 4781 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 7892 4781 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 7804 4781 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 7716 4781 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 7628 4781 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 7540 4781 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 7452 4781 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4741 7364 4781 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4728 10499 4792 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4728 10415 4792 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4728 10331 4792 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4661 7980 4701 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4661 7892 4701 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4661 7804 4701 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4661 7716 4701 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4661 7628 4701 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4661 7540 4701 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4661 7452 4701 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4661 7364 4701 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4660 11294 4700 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4660 9560 4700 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4647 10499 4711 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4647 10415 4711 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4647 10331 4711 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4581 7980 4621 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4581 7892 4621 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4581 7804 4621 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4581 7716 4621 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4581 7628 4621 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4581 7540 4621 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4581 7452 4621 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4581 7364 4621 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4579 11294 4619 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4579 9560 4619 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4566 10499 4630 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4566 10415 4630 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4566 10331 4630 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4501 7980 4541 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4501 7892 4541 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4501 7804 4541 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4501 7716 4541 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4501 7628 4541 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4501 7540 4541 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4501 7452 4541 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4501 7364 4541 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4498 11294 4538 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4498 9560 4538 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4485 10499 4549 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4485 10415 4549 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4485 10331 4549 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4421 7980 4461 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4421 7892 4461 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4421 7804 4461 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4421 7716 4461 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4421 7628 4461 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4421 7540 4461 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4421 7452 4461 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4421 7364 4461 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4417 11294 4457 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4417 9560 4457 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4404 10499 4468 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4404 10415 4468 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4404 10331 4468 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4341 7980 4381 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4341 7892 4381 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4341 7804 4381 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4341 7716 4381 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4341 7628 4381 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4341 7540 4381 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4341 7452 4381 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4341 7364 4381 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4336 11294 4376 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4336 9560 4376 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4323 10499 4387 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4323 10415 4387 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4323 10331 4387 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4261 7980 4301 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4261 7892 4301 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4261 7804 4301 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4261 7716 4301 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4261 7628 4301 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4261 7540 4301 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4261 7452 4301 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4261 7364 4301 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4255 11294 4295 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4255 9560 4295 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4242 10499 4306 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4242 10415 4306 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4242 10331 4306 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4181 7980 4221 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4181 7892 4221 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4181 7804 4221 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4181 7716 4221 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4181 7628 4221 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4181 7540 4221 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4181 7452 4221 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4181 7364 4221 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4174 11294 4214 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4174 9560 4214 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4161 10499 4225 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4161 10415 4225 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4161 10331 4225 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4100 7980 4140 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4100 7892 4140 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4100 7804 4140 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4100 7716 4140 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4100 7628 4140 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4100 7540 4140 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4100 7452 4140 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4100 7364 4140 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4093 11294 4133 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4093 9560 4133 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4080 10499 4144 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4080 10415 4144 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4080 10331 4144 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4019 7980 4059 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4019 7892 4059 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4019 7804 4059 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4019 7716 4059 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4019 7628 4059 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4019 7540 4059 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4019 7452 4059 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4019 7364 4059 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4012 11294 4052 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 4012 9560 4052 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3999 10499 4063 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3999 10415 4063 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3999 10331 4063 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3938 7980 3978 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3938 7892 3978 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3938 7804 3978 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3938 7716 3978 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3938 7628 3978 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3938 7540 3978 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3938 7452 3978 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3938 7364 3978 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3931 11294 3971 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3931 9560 3971 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3918 10499 3982 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3918 10415 3982 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3918 10331 3982 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3857 7980 3897 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3857 7892 3897 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3857 7804 3897 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3857 7716 3897 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3857 7628 3897 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3857 7540 3897 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3857 7452 3897 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3857 7364 3897 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3850 11294 3890 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3850 9560 3890 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3837 10499 3901 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3837 10415 3901 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3837 10331 3901 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3776 7980 3816 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3776 7892 3816 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3776 7804 3816 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3776 7716 3816 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3776 7628 3816 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3776 7540 3816 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3776 7452 3816 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3776 7364 3816 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3769 11294 3809 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3769 9560 3809 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3756 10499 3820 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3756 10415 3820 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3756 10331 3820 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3695 7980 3735 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3695 7892 3735 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3695 7804 3735 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3695 7716 3735 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3695 7628 3735 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3695 7540 3735 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3695 7452 3735 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3695 7364 3735 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3688 11294 3728 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3688 9560 3728 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3675 10499 3739 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3675 10415 3739 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3675 10331 3739 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3614 7980 3654 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3614 7892 3654 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3614 7804 3654 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3614 7716 3654 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3614 7628 3654 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3614 7540 3654 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3614 7452 3654 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3614 7364 3654 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3607 11294 3647 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3607 9560 3647 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3594 10499 3658 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3594 10415 3658 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3594 10331 3658 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3533 7980 3573 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3533 7892 3573 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3533 7804 3573 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3533 7716 3573 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3533 7628 3573 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3533 7540 3573 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3533 7452 3573 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3533 7364 3573 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3526 11294 3566 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3526 9560 3566 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3513 10499 3577 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3513 10415 3577 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3513 10331 3577 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3452 7980 3492 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3452 7892 3492 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3452 7804 3492 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3452 7716 3492 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3452 7628 3492 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3452 7540 3492 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3452 7452 3492 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3452 7364 3492 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3445 11294 3485 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3445 9560 3485 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3432 10499 3496 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3432 10415 3496 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3432 10331 3496 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3371 7980 3411 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3371 7892 3411 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3371 7804 3411 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3371 7716 3411 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3371 7628 3411 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3371 7540 3411 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3371 7452 3411 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3371 7364 3411 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3364 11294 3404 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3364 9560 3404 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3351 10499 3415 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3351 10415 3415 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3351 10331 3415 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3290 7980 3330 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3290 7892 3330 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3290 7804 3330 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3290 7716 3330 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3290 7628 3330 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3290 7540 3330 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3290 7452 3330 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3290 7364 3330 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3283 11294 3323 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3283 9560 3323 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3270 10499 3334 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3270 10415 3334 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3270 10331 3334 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3209 7980 3249 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3209 7892 3249 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3209 7804 3249 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3209 7716 3249 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3209 7628 3249 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3209 7540 3249 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3209 7452 3249 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3209 7364 3249 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3202 11294 3242 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3202 9560 3242 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3189 10499 3253 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3189 10415 3253 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3189 10331 3253 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3128 7980 3168 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3128 7892 3168 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3128 7804 3168 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3128 7716 3168 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3128 7628 3168 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3128 7540 3168 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3128 7452 3168 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3128 7364 3168 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3121 11294 3161 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3121 9560 3161 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3108 10499 3172 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3108 10415 3172 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3108 10331 3172 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3047 7980 3087 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3047 7892 3087 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3047 7804 3087 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3047 7716 3087 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3047 7628 3087 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3047 7540 3087 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3047 7452 3087 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3047 7364 3087 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3040 11294 3080 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3040 9560 3080 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3027 10499 3091 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3027 10415 3091 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 3027 10331 3091 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2966 7980 3006 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2966 7892 3006 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2966 7804 3006 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2966 7716 3006 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2966 7628 3006 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2966 7540 3006 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2966 7452 3006 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2966 7364 3006 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2959 11294 2999 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2959 9560 2999 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2946 10499 3010 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2946 10415 3010 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2946 10331 3010 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2885 7980 2925 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2885 7892 2925 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2885 7804 2925 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2885 7716 2925 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2885 7628 2925 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2885 7540 2925 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2885 7452 2925 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2885 7364 2925 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2878 11294 2918 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2878 9560 2918 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2865 10499 2929 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2865 10415 2929 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2865 10331 2929 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2804 7980 2844 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2804 7892 2844 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2804 7804 2844 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2804 7716 2844 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2804 7628 2844 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2804 7540 2844 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2804 7452 2844 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2804 7364 2844 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2797 11294 2837 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2797 9560 2837 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2784 10499 2848 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2784 10415 2848 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2784 10331 2848 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2723 7980 2763 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2723 7892 2763 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2723 7804 2763 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2723 7716 2763 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2723 7628 2763 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2723 7540 2763 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2723 7452 2763 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2723 7364 2763 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2716 11294 2756 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2716 9560 2756 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2703 10499 2767 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2703 10415 2767 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2703 10331 2767 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2642 7980 2682 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2642 7892 2682 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2642 7804 2682 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2642 7716 2682 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2642 7628 2682 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2642 7540 2682 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2642 7452 2682 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2642 7364 2682 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2635 11294 2675 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2635 9560 2675 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2622 10499 2686 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2622 10415 2686 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2622 10331 2686 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2561 7980 2601 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2561 7892 2601 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2561 7804 2601 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2561 7716 2601 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2561 7628 2601 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2561 7540 2601 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2561 7452 2601 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2561 7364 2601 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2554 11294 2594 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2554 9560 2594 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2541 10499 2605 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2541 10415 2605 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2541 10331 2605 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2480 7980 2520 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2480 7892 2520 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2480 7804 2520 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2480 7716 2520 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2480 7628 2520 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2480 7540 2520 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2480 7452 2520 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2480 7364 2520 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2473 11294 2513 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2473 9560 2513 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2460 10499 2524 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2460 10415 2524 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2460 10331 2524 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2399 7980 2439 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2399 7892 2439 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2399 7804 2439 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2399 7716 2439 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2399 7628 2439 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2399 7540 2439 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2399 7452 2439 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2399 7364 2439 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2392 11294 2432 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2392 9560 2432 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2379 10499 2443 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2379 10415 2443 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2379 10331 2443 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2318 7980 2358 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2318 7892 2358 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2318 7804 2358 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2318 7716 2358 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2318 7628 2358 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2318 7540 2358 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2318 7452 2358 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2318 7364 2358 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2311 11294 2351 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2311 9560 2351 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2298 10499 2362 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2298 10415 2362 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2298 10331 2362 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2237 7980 2277 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2237 7892 2277 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2237 7804 2277 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2237 7716 2277 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2237 7628 2277 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2237 7540 2277 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2237 7452 2277 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2237 7364 2277 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2230 11294 2270 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2230 9560 2270 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2217 10499 2281 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2217 10415 2281 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2217 10331 2281 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2156 7980 2196 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2156 7892 2196 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2156 7804 2196 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2156 7716 2196 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2156 7628 2196 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2156 7540 2196 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2156 7452 2196 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2156 7364 2196 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2149 11294 2189 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2149 9560 2189 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2136 10499 2200 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2136 10415 2200 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2136 10331 2200 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2075 7980 2115 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2075 7892 2115 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2075 7804 2115 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2075 7716 2115 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2075 7628 2115 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2075 7540 2115 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2075 7452 2115 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2075 7364 2115 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2068 11294 2108 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2068 9560 2108 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2055 10499 2119 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2055 10415 2119 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 2055 10331 2119 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1994 7980 2034 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1994 7892 2034 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1994 7804 2034 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1994 7716 2034 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1994 7628 2034 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1994 7540 2034 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1994 7452 2034 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1994 7364 2034 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1987 11294 2027 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1987 9560 2027 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1974 10499 2038 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1974 10415 2038 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1974 10331 2038 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1913 7980 1953 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1913 7892 1953 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1913 7804 1953 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1913 7716 1953 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1913 7628 1953 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1913 7540 1953 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1913 7452 1953 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1913 7364 1953 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1906 11294 1946 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1906 9560 1946 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1893 10499 1957 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1893 10415 1957 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1893 10331 1957 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1832 7980 1872 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1832 7892 1872 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1832 7804 1872 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1832 7716 1872 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1832 7628 1872 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1832 7540 1872 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1832 7452 1872 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1832 7364 1872 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1825 11294 1865 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1825 9560 1865 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1812 10499 1876 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1812 10415 1876 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1812 10331 1876 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1751 7980 1791 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1751 7892 1791 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1751 7804 1791 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1751 7716 1791 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1751 7628 1791 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1751 7540 1791 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1751 7452 1791 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1751 7364 1791 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1744 11294 1784 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1744 9560 1784 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1731 10499 1795 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1731 10415 1795 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1731 10331 1795 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1670 7980 1710 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1670 7892 1710 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1670 7804 1710 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1670 7716 1710 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1670 7628 1710 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1670 7540 1710 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1670 7452 1710 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1670 7364 1710 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1663 11294 1703 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1663 9560 1703 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1650 10499 1714 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1650 10415 1714 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1650 10331 1714 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1589 7980 1629 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1589 7892 1629 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1589 7804 1629 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1589 7716 1629 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1589 7628 1629 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1589 7540 1629 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1589 7452 1629 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1589 7364 1629 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1582 11294 1622 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1582 9560 1622 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1569 10499 1633 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1569 10415 1633 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1569 10331 1633 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1508 7980 1548 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1508 7892 1548 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1508 7804 1548 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1508 7716 1548 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1508 7628 1548 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1508 7540 1548 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1508 7452 1548 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1508 7364 1548 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1501 11294 1541 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1501 9560 1541 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1488 10499 1552 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1488 10415 1552 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1488 10331 1552 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1427 7980 1467 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1427 7892 1467 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1427 7804 1467 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1427 7716 1467 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1427 7628 1467 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1427 7540 1467 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1427 7452 1467 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1427 7364 1467 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1420 11294 1460 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1420 9560 1460 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1407 10499 1471 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1407 10415 1471 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1407 10331 1471 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1346 7980 1386 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1346 7892 1386 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1346 7804 1386 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1346 7716 1386 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1346 7628 1386 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1346 7540 1386 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1346 7452 1386 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1346 7364 1386 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1339 11294 1379 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1339 9560 1379 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1326 10499 1390 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1326 10415 1390 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1326 10331 1390 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1265 7980 1305 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1265 7892 1305 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1265 7804 1305 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1265 7716 1305 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1265 7628 1305 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1265 7540 1305 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1265 7452 1305 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1265 7364 1305 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1258 11294 1298 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1258 9560 1298 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1245 10499 1309 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1245 10415 1309 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1245 10331 1309 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1184 7980 1224 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1184 7892 1224 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1184 7804 1224 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1184 7716 1224 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1184 7628 1224 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1184 7540 1224 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1184 7452 1224 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1184 7364 1224 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1177 11294 1217 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1177 9560 1217 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1164 10499 1228 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1164 10415 1228 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1164 10331 1228 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1103 7980 1143 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1103 7892 1143 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1103 7804 1143 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1103 7716 1143 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1103 7628 1143 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1103 7540 1143 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1103 7452 1143 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1103 7364 1143 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1096 11294 1136 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1096 9560 1136 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1083 10499 1147 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1083 10415 1147 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1083 10331 1147 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1022 7980 1062 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1022 7892 1062 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1022 7804 1062 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1022 7716 1062 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1022 7628 1062 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1022 7540 1062 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1022 7452 1062 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1022 7364 1062 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1015 11294 1055 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1015 9560 1055 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1002 10499 1066 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1002 10415 1066 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 1002 10331 1066 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 941 7980 981 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 941 7892 981 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 941 7804 981 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 941 7716 981 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 941 7628 981 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 941 7540 981 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 941 7452 981 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 941 7364 981 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 934 11294 974 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 934 9560 974 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 921 10499 985 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 921 10415 985 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 921 10331 985 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 860 7980 900 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 860 7892 900 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 860 7804 900 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 860 7716 900 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 860 7628 900 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 860 7540 900 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 860 7452 900 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 860 7364 900 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 853 11294 893 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 853 9560 893 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 840 10499 904 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 840 10415 904 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 840 10331 904 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 779 7980 819 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 779 7892 819 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 779 7804 819 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 779 7716 819 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 779 7628 819 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 779 7540 819 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 779 7452 819 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 779 7364 819 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 772 11294 812 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 772 9560 812 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 759 10499 823 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 759 10415 823 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 759 10331 823 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 698 7980 738 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 698 7892 738 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 698 7804 738 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 698 7716 738 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 698 7628 738 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 698 7540 738 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 698 7452 738 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 698 7364 738 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 691 11294 731 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 691 9560 731 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 678 10499 742 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 678 10415 742 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 678 10331 742 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 617 7980 657 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 617 7892 657 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 617 7804 657 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 617 7716 657 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 617 7628 657 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 617 7540 657 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 617 7452 657 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 617 7364 657 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 610 11294 650 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 610 9560 650 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 597 10499 661 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 597 10415 661 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 597 10331 661 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 536 7980 576 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 536 7892 576 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 536 7804 576 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 536 7716 576 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 536 7628 576 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 536 7540 576 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 536 7452 576 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 536 7364 576 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 529 11294 569 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 529 9560 569 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 515 10499 579 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 515 10415 579 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 515 10331 579 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 455 7980 495 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 455 7892 495 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 455 7804 495 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 455 7716 495 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 455 7628 495 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 455 7540 495 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 455 7452 495 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 455 7364 495 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 448 11294 488 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 448 9560 488 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 433 10499 497 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 433 10415 497 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 433 10331 497 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 374 7980 414 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 374 7892 414 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 374 7804 414 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 374 7716 414 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 374 7628 414 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 374 7540 414 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 374 7452 414 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 374 7364 414 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 367 11294 407 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 367 9560 407 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 351 10499 415 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 351 10415 415 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 351 10331 415 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 293 7980 333 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 293 7892 333 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 293 7804 333 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 293 7716 333 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 293 7628 333 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 293 7540 333 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 293 7452 333 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 293 7364 333 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 286 11294 326 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 286 9560 326 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 269 10499 333 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 269 10415 333 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 269 10331 333 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 212 7980 252 8020 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 212 7892 252 7932 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 212 7804 252 7844 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 212 7716 252 7756 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 212 7628 252 7668 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 212 7540 252 7580 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 212 7452 252 7492 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 212 7364 252 7404 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 205 11294 245 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 205 9560 245 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 187 10499 251 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 187 10415 251 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 187 10331 251 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 124 11294 164 11334 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 124 9560 164 9600 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 105 10499 169 10563 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 105 10415 169 10479 6 VSSA
port 40 nsew ground bidirectional
rlabel metal3 s 105 10331 169 10395 6 VSSA
port 40 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 41 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 42 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 43 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 44 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 44 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 44 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 44 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 45 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 46 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 47 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 48 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 49 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 50 nsew ground bidirectional
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 52 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 53 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 54 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 56 nsew ground bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 57 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 58 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 59 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 60 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 60 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 60 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 60 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 25819050
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25712154
<< end >>
