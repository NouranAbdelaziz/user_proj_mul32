/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/klayout/pymacros/cells/fixed_devices/VPP/sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield.cdl