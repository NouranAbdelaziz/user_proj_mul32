magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal4 >>
rect 0 35890 287 40733
rect 0 14740 529 19733
rect 0 13550 296 14440
rect 0 12380 325 13270
rect 0 11358 4582 11954
rect 0 10406 4187 11002
rect 0 9050 295 9980
rect 0 7110 277 7800
rect 0 5900 320 6830
rect 0 4690 305 5620
rect 0 3720 294 4410
rect 0 2510 757 3440
rect 0 1140 470 2230
rect 407 0 1497 254
rect 1777 0 2707 254
rect 2987 0 3677 251
rect 3957 0 4887 254
rect 6377 0 7067 254
rect 8317 0 9247 254
rect 9673 0 10269 4175
rect 10625 0 11221 3695
rect 11647 0 12537 254
rect 12817 0 13707 254
rect 14007 0 19000 304
<< obsm4 >>
rect 367 35810 40000 40733
rect 0 19813 40000 35810
rect 609 14660 40000 19813
rect 0 14520 40000 14660
rect 376 13470 40000 14520
rect 0 13350 40000 13470
rect 405 12300 40000 13350
rect 0 12034 40000 12300
rect 0 12014 4635 12034
rect 0 11278 4310 11298
rect 4662 11278 40000 12034
rect 0 11062 40000 11278
rect 0 10326 3915 10346
rect 4267 10326 40000 11062
rect 0 10060 40000 10326
rect 375 8970 40000 10060
rect 0 7880 40000 8970
rect 357 7030 40000 7880
rect 0 6910 40000 7030
rect 400 5820 40000 6910
rect 0 5700 40000 5820
rect 385 4610 40000 5700
rect 0 4490 40000 4610
rect 374 4255 40000 4490
rect 374 3640 9593 4255
rect 0 3520 9593 3640
rect 837 2430 9593 3520
rect 0 2310 9593 2430
tri 0 1060 80 1140 ne
rect 80 1060 407 1140
rect 550 1060 9593 2310
rect 0 334 9593 1060
rect 0 0 327 334
rect 1577 0 1697 334
rect 2787 331 3877 334
rect 2787 0 2907 331
rect 3757 0 3877 331
rect 4967 0 6297 334
rect 7147 0 8237 334
rect 9327 0 9593 334
rect 10349 3775 40000 4255
rect 10349 0 10545 3775
rect 11301 384 40000 3775
rect 11301 334 13927 384
rect 11301 0 11567 334
rect 12617 0 12737 334
rect 13787 0 13927 334
rect 19080 0 40000 384
<< metal5 >>
rect 0 35890 287 40733
rect 0 14740 529 19730
rect 0 13570 296 14420
rect 0 12400 325 13250
rect 0 10280 4631 12080
rect 0 9070 295 9960
rect 0 7130 277 7780
rect 0 5920 320 6810
rect 0 4710 305 5600
rect 0 3740 294 4390
rect 0 2530 757 3420
rect 0 1160 470 2210
rect 427 0 1477 254
rect 1797 0 2687 254
rect 3007 0 3657 251
rect 3977 0 4867 254
rect 5187 0 6077 254
rect 6397 0 7047 254
rect 8337 0 9227 254
rect 11667 0 12517 254
rect 12837 0 13687 254
rect 14007 0 18997 304
rect 35157 0 40000 254
<< obsm5 >>
rect 607 35570 40000 40733
rect 0 20050 40000 35570
rect 849 14420 40000 20050
rect 616 13570 40000 14420
rect 645 12400 40000 13570
rect 4951 9960 40000 12400
rect 615 8750 40000 9960
rect 0 8100 40000 8750
rect 597 7130 40000 8100
rect 640 5600 40000 7130
rect 625 4390 40000 5600
rect 614 3740 40000 4390
rect 1077 2210 40000 3740
tri 0 840 320 1160 ne
rect 320 840 427 1160
rect 790 840 40000 2210
rect 0 624 40000 840
rect 0 574 13687 624
rect 19317 574 40000 624
rect 0 0 107 574
rect 3007 571 3657 574
rect 7367 0 8017 574
rect 9547 0 11347 574
rect 19317 0 34837 574
<< labels >>
rlabel metal4 s 0 11358 4582 11954 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 10625 0 11221 3695 6 AMUXBUS_A
port 2 nsew signal bidirectional
rlabel metal4 s 0 10406 4187 11002 6 AMUXBUS_B
port 3 nsew signal bidirectional
rlabel metal4 s 9673 0 10269 4175 6 AMUXBUS_B
port 4 nsew signal bidirectional
rlabel metal5 s 0 2530 757 3420 6 VCCD
port 5 nsew signal bidirectional
rlabel metal5 s 1797 0 2687 254 6 VCCD
port 6 nsew signal bidirectional
rlabel metal4 s 0 2510 757 3440 6 VCCD
port 7 nsew signal bidirectional
rlabel metal4 s 1777 0 2707 254 6 VCCD
port 8 nsew signal bidirectional
rlabel metal5 s 0 1160 470 2210 6 VCCHIB
port 9 nsew signal bidirectional
rlabel metal5 s 427 0 1477 254 6 VCCHIB
port 10 nsew signal bidirectional
rlabel metal4 s 0 1140 470 2230 6 VCCHIB
port 11 nsew signal bidirectional
rlabel metal4 s 407 0 1497 254 6 VCCHIB
port 12 nsew signal bidirectional
rlabel metal5 s 0 3740 294 4390 6 VDDA
port 13 nsew signal bidirectional
rlabel metal5 s 3007 0 3657 251 6 VDDA
port 14 nsew signal bidirectional
rlabel metal4 s 0 3720 294 4410 6 VDDA
port 15 nsew signal bidirectional
rlabel metal4 s 2987 0 3677 251 6 VDDA
port 16 nsew signal bidirectional
rlabel metal5 s 0 14740 529 19730 6 VDDIO
port 17 nsew signal bidirectional
rlabel metal5 s 0 4710 305 5600 6 VDDIO
port 18 nsew signal bidirectional
rlabel metal5 s 3977 0 4867 254 6 VDDIO
port 19 nsew signal bidirectional
rlabel metal5 s 14007 0 18997 304 6 VDDIO
port 20 nsew signal bidirectional
rlabel metal4 s 0 4690 305 5620 6 VDDIO
port 21 nsew signal bidirectional
rlabel metal4 s 0 14740 529 19733 6 VDDIO
port 22 nsew signal bidirectional
rlabel metal4 s 14007 0 19000 304 6 VDDIO
port 23 nsew signal bidirectional
rlabel metal4 s 3957 0 4887 254 6 VDDIO
port 24 nsew signal bidirectional
rlabel metal5 s 0 13570 296 14420 6 VDDIO_Q
port 25 nsew signal bidirectional
rlabel metal5 s 12837 0 13687 254 6 VDDIO_Q
port 26 nsew signal bidirectional
rlabel metal4 s 0 13550 296 14440 6 VDDIO_Q
port 27 nsew signal bidirectional
rlabel metal4 s 12817 0 13707 254 6 VDDIO_Q
port 28 nsew signal bidirectional
rlabel metal5 s 0 10280 4631 12080 6 VSSA
port 29 nsew signal bidirectional
rlabel metal5 s 0 9070 295 9960 6 VSSD
port 30 nsew signal bidirectional
rlabel metal5 s 8337 0 9227 254 6 VSSD
port 31 nsew signal bidirectional
rlabel metal4 s 0 9050 295 9980 6 VSSD
port 32 nsew signal bidirectional
rlabel metal4 s 8317 0 9247 254 6 VSSD
port 33 nsew signal bidirectional
rlabel metal5 s 0 35890 287 40733 6 VSSIO
port 34 nsew signal bidirectional
rlabel metal5 s 0 5920 320 6810 6 VSSIO
port 35 nsew signal bidirectional
rlabel metal5 s 5187 0 6077 254 6 VSSIO
port 36 nsew signal bidirectional
rlabel metal5 s 35157 0 40000 254 6 VSSIO
port 37 nsew signal bidirectional
rlabel metal4 s 0 5900 320 6830 6 VSSIO
port 38 nsew signal bidirectional
rlabel metal4 s 0 35890 287 40733 6 VSSIO
port 39 nsew signal bidirectional
rlabel metal5 s 0 12400 325 13250 6 VSSIO_Q
port 40 nsew signal bidirectional
rlabel metal5 s 11667 0 12517 254 6 VSSIO_Q
port 41 nsew signal bidirectional
rlabel metal4 s 0 12380 325 13270 6 VSSIO_Q
port 42 nsew signal bidirectional
rlabel metal4 s 11647 0 12537 254 6 VSSIO_Q
port 43 nsew signal bidirectional
rlabel metal5 s 0 7130 277 7780 6 VSWITCH
port 44 nsew signal bidirectional
rlabel metal5 s 6397 0 7047 254 6 VSWITCH
port 45 nsew signal bidirectional
rlabel metal4 s 0 7110 277 7800 6 VSWITCH
port 46 nsew signal bidirectional
rlabel metal4 s 6377 0 7067 254 6 VSWITCH
port 47 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40733
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 27794742
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27529686
<< end >>
