magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal3 >>
rect 99 39983 14858 40000
rect 99 39919 125 39983
rect 189 39919 205 39983
rect 269 39919 285 39983
rect 349 39919 365 39983
rect 429 39919 445 39983
rect 509 39919 525 39983
rect 589 39919 605 39983
rect 669 39919 685 39983
rect 749 39919 765 39983
rect 829 39919 845 39983
rect 909 39919 925 39983
rect 989 39919 1005 39983
rect 1069 39919 1085 39983
rect 1149 39919 1165 39983
rect 1229 39919 1245 39983
rect 1309 39919 1325 39983
rect 1389 39919 1405 39983
rect 1469 39919 1485 39983
rect 1549 39919 1565 39983
rect 1629 39919 1645 39983
rect 1709 39919 1725 39983
rect 1789 39919 1805 39983
rect 1869 39919 1885 39983
rect 1949 39919 1965 39983
rect 2029 39919 2045 39983
rect 2109 39919 2125 39983
rect 2189 39919 2205 39983
rect 2269 39919 2285 39983
rect 2349 39919 2365 39983
rect 2429 39919 2445 39983
rect 2509 39919 2525 39983
rect 2589 39919 2605 39983
rect 2669 39982 12306 39983
rect 2669 39919 2727 39982
rect 99 39918 2727 39919
rect 2791 39918 2808 39982
rect 2872 39918 2889 39982
rect 2953 39918 2970 39982
rect 3034 39918 3051 39982
rect 3115 39918 3132 39982
rect 3196 39918 3213 39982
rect 3277 39918 3294 39982
rect 3358 39918 3375 39982
rect 3439 39918 3456 39982
rect 3520 39918 3537 39982
rect 3601 39918 3618 39982
rect 3682 39918 3699 39982
rect 3763 39918 3780 39982
rect 3844 39918 3861 39982
rect 3925 39918 3942 39982
rect 4006 39918 4023 39982
rect 4087 39918 4104 39982
rect 4168 39918 4185 39982
rect 4249 39918 4266 39982
rect 4330 39918 4347 39982
rect 4411 39918 4428 39982
rect 4492 39918 4509 39982
rect 4573 39918 4590 39982
rect 4654 39918 4671 39982
rect 4735 39918 4752 39982
rect 4816 39918 4833 39982
rect 4897 39918 4914 39982
rect 4978 39918 4995 39982
rect 5059 39918 5076 39982
rect 5140 39918 5157 39982
rect 5221 39918 5238 39982
rect 5302 39918 5319 39982
rect 5383 39918 5400 39982
rect 99 39902 5400 39918
rect 99 39838 125 39902
rect 189 39838 205 39902
rect 269 39838 285 39902
rect 349 39838 365 39902
rect 429 39838 445 39902
rect 509 39838 525 39902
rect 589 39838 605 39902
rect 669 39838 685 39902
rect 749 39838 765 39902
rect 829 39838 845 39902
rect 909 39838 925 39902
rect 989 39838 1005 39902
rect 1069 39838 1085 39902
rect 1149 39838 1165 39902
rect 1229 39838 1245 39902
rect 1309 39838 1325 39902
rect 1389 39838 1405 39902
rect 1469 39838 1485 39902
rect 1549 39838 1565 39902
rect 1629 39838 1645 39902
rect 1709 39838 1725 39902
rect 1789 39838 1805 39902
rect 1869 39838 1885 39902
rect 1949 39838 1965 39902
rect 2029 39838 2045 39902
rect 2109 39838 2125 39902
rect 2189 39838 2205 39902
rect 2269 39838 2285 39902
rect 2349 39838 2365 39902
rect 2429 39838 2445 39902
rect 2509 39838 2525 39902
rect 2589 39838 2605 39902
rect 2669 39838 2727 39902
rect 2791 39838 2808 39902
rect 2872 39838 2889 39902
rect 2953 39838 2970 39902
rect 3034 39838 3051 39902
rect 3115 39838 3132 39902
rect 3196 39838 3213 39902
rect 3277 39838 3294 39902
rect 3358 39838 3375 39902
rect 3439 39838 3456 39902
rect 3520 39838 3537 39902
rect 3601 39838 3618 39902
rect 3682 39838 3699 39902
rect 3763 39838 3780 39902
rect 3844 39838 3861 39902
rect 3925 39838 3942 39902
rect 4006 39838 4023 39902
rect 4087 39838 4104 39902
rect 4168 39838 4185 39902
rect 4249 39838 4266 39902
rect 4330 39838 4347 39902
rect 4411 39838 4428 39902
rect 4492 39838 4509 39902
rect 4573 39838 4590 39902
rect 4654 39838 4671 39902
rect 4735 39838 4752 39902
rect 4816 39838 4833 39902
rect 4897 39838 4914 39902
rect 4978 39838 4995 39902
rect 5059 39838 5076 39902
rect 5140 39838 5157 39902
rect 5221 39838 5238 39902
rect 5302 39838 5319 39902
rect 5383 39838 5400 39902
rect 99 39822 5400 39838
rect 99 39821 2727 39822
rect 99 39757 125 39821
rect 189 39757 205 39821
rect 269 39757 285 39821
rect 349 39757 365 39821
rect 429 39757 445 39821
rect 509 39757 525 39821
rect 589 39757 605 39821
rect 669 39757 685 39821
rect 749 39757 765 39821
rect 829 39757 845 39821
rect 909 39757 925 39821
rect 989 39757 1005 39821
rect 1069 39757 1085 39821
rect 1149 39757 1165 39821
rect 1229 39757 1245 39821
rect 1309 39757 1325 39821
rect 1389 39757 1405 39821
rect 1469 39757 1485 39821
rect 1549 39757 1565 39821
rect 1629 39757 1645 39821
rect 1709 39757 1725 39821
rect 1789 39757 1805 39821
rect 1869 39757 1885 39821
rect 1949 39757 1965 39821
rect 2029 39757 2045 39821
rect 2109 39757 2125 39821
rect 2189 39757 2205 39821
rect 2269 39757 2285 39821
rect 2349 39757 2365 39821
rect 2429 39757 2445 39821
rect 2509 39757 2525 39821
rect 2589 39757 2605 39821
rect 2669 39758 2727 39821
rect 2791 39758 2808 39822
rect 2872 39758 2889 39822
rect 2953 39758 2970 39822
rect 3034 39758 3051 39822
rect 3115 39758 3132 39822
rect 3196 39758 3213 39822
rect 3277 39758 3294 39822
rect 3358 39758 3375 39822
rect 3439 39758 3456 39822
rect 3520 39758 3537 39822
rect 3601 39758 3618 39822
rect 3682 39758 3699 39822
rect 3763 39758 3780 39822
rect 3844 39758 3861 39822
rect 3925 39758 3942 39822
rect 4006 39758 4023 39822
rect 4087 39758 4104 39822
rect 4168 39758 4185 39822
rect 4249 39758 4266 39822
rect 4330 39758 4347 39822
rect 4411 39758 4428 39822
rect 4492 39758 4509 39822
rect 4573 39758 4590 39822
rect 4654 39758 4671 39822
rect 4735 39758 4752 39822
rect 4816 39758 4833 39822
rect 4897 39758 4914 39822
rect 4978 39758 4995 39822
rect 5059 39758 5076 39822
rect 5140 39758 5157 39822
rect 5221 39758 5238 39822
rect 5302 39758 5319 39822
rect 5383 39758 5400 39822
rect 2669 39757 5400 39758
rect 99 39742 5400 39757
rect 99 39740 2727 39742
rect 99 39676 125 39740
rect 189 39676 205 39740
rect 269 39676 285 39740
rect 349 39676 365 39740
rect 429 39676 445 39740
rect 509 39676 525 39740
rect 589 39676 605 39740
rect 669 39676 685 39740
rect 749 39676 765 39740
rect 829 39676 845 39740
rect 909 39676 925 39740
rect 989 39676 1005 39740
rect 1069 39676 1085 39740
rect 1149 39676 1165 39740
rect 1229 39676 1245 39740
rect 1309 39676 1325 39740
rect 1389 39676 1405 39740
rect 1469 39676 1485 39740
rect 1549 39676 1565 39740
rect 1629 39676 1645 39740
rect 1709 39676 1725 39740
rect 1789 39676 1805 39740
rect 1869 39676 1885 39740
rect 1949 39676 1965 39740
rect 2029 39676 2045 39740
rect 2109 39676 2125 39740
rect 2189 39676 2205 39740
rect 2269 39676 2285 39740
rect 2349 39676 2365 39740
rect 2429 39676 2445 39740
rect 2509 39676 2525 39740
rect 2589 39676 2605 39740
rect 2669 39678 2727 39740
rect 2791 39678 2808 39742
rect 2872 39678 2889 39742
rect 2953 39678 2970 39742
rect 3034 39678 3051 39742
rect 3115 39678 3132 39742
rect 3196 39678 3213 39742
rect 3277 39678 3294 39742
rect 3358 39678 3375 39742
rect 3439 39678 3456 39742
rect 3520 39678 3537 39742
rect 3601 39678 3618 39742
rect 3682 39678 3699 39742
rect 3763 39678 3780 39742
rect 3844 39678 3861 39742
rect 3925 39678 3942 39742
rect 4006 39678 4023 39742
rect 4087 39678 4104 39742
rect 4168 39678 4185 39742
rect 4249 39678 4266 39742
rect 4330 39678 4347 39742
rect 4411 39678 4428 39742
rect 4492 39678 4509 39742
rect 4573 39678 4590 39742
rect 4654 39678 4671 39742
rect 4735 39678 4752 39742
rect 4816 39678 4833 39742
rect 4897 39678 4914 39742
rect 4978 39678 4995 39742
rect 5059 39678 5076 39742
rect 5140 39678 5157 39742
rect 5221 39678 5238 39742
rect 5302 39678 5319 39742
rect 5383 39678 5400 39742
rect 2669 39676 5400 39678
rect 99 39662 5400 39676
rect 99 39659 2727 39662
rect 99 39595 125 39659
rect 189 39595 205 39659
rect 269 39595 285 39659
rect 349 39595 365 39659
rect 429 39595 445 39659
rect 509 39595 525 39659
rect 589 39595 605 39659
rect 669 39595 685 39659
rect 749 39595 765 39659
rect 829 39595 845 39659
rect 909 39595 925 39659
rect 989 39595 1005 39659
rect 1069 39595 1085 39659
rect 1149 39595 1165 39659
rect 1229 39595 1245 39659
rect 1309 39595 1325 39659
rect 1389 39595 1405 39659
rect 1469 39595 1485 39659
rect 1549 39595 1565 39659
rect 1629 39595 1645 39659
rect 1709 39595 1725 39659
rect 1789 39595 1805 39659
rect 1869 39595 1885 39659
rect 1949 39595 1965 39659
rect 2029 39595 2045 39659
rect 2109 39595 2125 39659
rect 2189 39595 2205 39659
rect 2269 39595 2285 39659
rect 2349 39595 2365 39659
rect 2429 39595 2445 39659
rect 2509 39595 2525 39659
rect 2589 39595 2605 39659
rect 2669 39598 2727 39659
rect 2791 39598 2808 39662
rect 2872 39598 2889 39662
rect 2953 39598 2970 39662
rect 3034 39598 3051 39662
rect 3115 39598 3132 39662
rect 3196 39598 3213 39662
rect 3277 39598 3294 39662
rect 3358 39598 3375 39662
rect 3439 39598 3456 39662
rect 3520 39598 3537 39662
rect 3601 39598 3618 39662
rect 3682 39598 3699 39662
rect 3763 39598 3780 39662
rect 3844 39598 3861 39662
rect 3925 39598 3942 39662
rect 4006 39598 4023 39662
rect 4087 39598 4104 39662
rect 4168 39598 4185 39662
rect 4249 39598 4266 39662
rect 4330 39598 4347 39662
rect 4411 39598 4428 39662
rect 4492 39598 4509 39662
rect 4573 39598 4590 39662
rect 4654 39598 4671 39662
rect 4735 39598 4752 39662
rect 4816 39598 4833 39662
rect 4897 39598 4914 39662
rect 4978 39598 4995 39662
rect 5059 39598 5076 39662
rect 5140 39598 5157 39662
rect 5221 39598 5238 39662
rect 5302 39598 5319 39662
rect 5383 39598 5400 39662
rect 2669 39595 5400 39598
rect 99 39582 5400 39595
rect 99 39578 2727 39582
rect 99 39514 125 39578
rect 189 39514 205 39578
rect 269 39514 285 39578
rect 349 39514 365 39578
rect 429 39514 445 39578
rect 509 39514 525 39578
rect 589 39514 605 39578
rect 669 39514 685 39578
rect 749 39514 765 39578
rect 829 39514 845 39578
rect 909 39514 925 39578
rect 989 39514 1005 39578
rect 1069 39514 1085 39578
rect 1149 39514 1165 39578
rect 1229 39514 1245 39578
rect 1309 39514 1325 39578
rect 1389 39514 1405 39578
rect 1469 39514 1485 39578
rect 1549 39514 1565 39578
rect 1629 39514 1645 39578
rect 1709 39514 1725 39578
rect 1789 39514 1805 39578
rect 1869 39514 1885 39578
rect 1949 39514 1965 39578
rect 2029 39514 2045 39578
rect 2109 39514 2125 39578
rect 2189 39514 2205 39578
rect 2269 39514 2285 39578
rect 2349 39514 2365 39578
rect 2429 39514 2445 39578
rect 2509 39514 2525 39578
rect 2589 39514 2605 39578
rect 2669 39518 2727 39578
rect 2791 39518 2808 39582
rect 2872 39518 2889 39582
rect 2953 39518 2970 39582
rect 3034 39518 3051 39582
rect 3115 39518 3132 39582
rect 3196 39518 3213 39582
rect 3277 39518 3294 39582
rect 3358 39518 3375 39582
rect 3439 39518 3456 39582
rect 3520 39518 3537 39582
rect 3601 39518 3618 39582
rect 3682 39518 3699 39582
rect 3763 39518 3780 39582
rect 3844 39518 3861 39582
rect 3925 39518 3942 39582
rect 4006 39518 4023 39582
rect 4087 39518 4104 39582
rect 4168 39518 4185 39582
rect 4249 39518 4266 39582
rect 4330 39518 4347 39582
rect 4411 39518 4428 39582
rect 4492 39518 4509 39582
rect 4573 39518 4590 39582
rect 4654 39518 4671 39582
rect 4735 39518 4752 39582
rect 4816 39518 4833 39582
rect 4897 39518 4914 39582
rect 4978 39518 4995 39582
rect 5059 39518 5076 39582
rect 5140 39518 5157 39582
rect 5221 39518 5238 39582
rect 5302 39518 5319 39582
rect 5383 39518 5400 39582
rect 2669 39514 5400 39518
rect 99 39502 5400 39514
rect 99 39497 2727 39502
rect 99 39433 125 39497
rect 189 39433 205 39497
rect 269 39433 285 39497
rect 349 39433 365 39497
rect 429 39433 445 39497
rect 509 39433 525 39497
rect 589 39433 605 39497
rect 669 39433 685 39497
rect 749 39433 765 39497
rect 829 39433 845 39497
rect 909 39433 925 39497
rect 989 39433 1005 39497
rect 1069 39433 1085 39497
rect 1149 39433 1165 39497
rect 1229 39433 1245 39497
rect 1309 39433 1325 39497
rect 1389 39433 1405 39497
rect 1469 39433 1485 39497
rect 1549 39433 1565 39497
rect 1629 39433 1645 39497
rect 1709 39433 1725 39497
rect 1789 39433 1805 39497
rect 1869 39433 1885 39497
rect 1949 39433 1965 39497
rect 2029 39433 2045 39497
rect 2109 39433 2125 39497
rect 2189 39433 2205 39497
rect 2269 39433 2285 39497
rect 2349 39433 2365 39497
rect 2429 39433 2445 39497
rect 2509 39433 2525 39497
rect 2589 39433 2605 39497
rect 2669 39438 2727 39497
rect 2791 39438 2808 39502
rect 2872 39438 2889 39502
rect 2953 39438 2970 39502
rect 3034 39438 3051 39502
rect 3115 39438 3132 39502
rect 3196 39438 3213 39502
rect 3277 39438 3294 39502
rect 3358 39438 3375 39502
rect 3439 39438 3456 39502
rect 3520 39438 3537 39502
rect 3601 39438 3618 39502
rect 3682 39438 3699 39502
rect 3763 39438 3780 39502
rect 3844 39438 3861 39502
rect 3925 39438 3942 39502
rect 4006 39438 4023 39502
rect 4087 39438 4104 39502
rect 4168 39438 4185 39502
rect 4249 39438 4266 39502
rect 4330 39438 4347 39502
rect 4411 39438 4428 39502
rect 4492 39438 4509 39502
rect 4573 39438 4590 39502
rect 4654 39438 4671 39502
rect 4735 39438 4752 39502
rect 4816 39438 4833 39502
rect 4897 39438 4914 39502
rect 4978 39438 4995 39502
rect 5059 39438 5076 39502
rect 5140 39438 5157 39502
rect 5221 39438 5238 39502
rect 5302 39438 5319 39502
rect 5383 39438 5400 39502
rect 12264 39919 12306 39982
rect 12370 39919 12386 39983
rect 12450 39919 12466 39983
rect 12530 39919 12546 39983
rect 12610 39919 12626 39983
rect 12690 39919 12706 39983
rect 12770 39919 12786 39983
rect 12850 39919 12866 39983
rect 12930 39919 12946 39983
rect 13010 39919 13026 39983
rect 13090 39919 13106 39983
rect 13170 39919 13186 39983
rect 13250 39919 13266 39983
rect 13330 39919 13346 39983
rect 13410 39919 13426 39983
rect 13490 39919 13506 39983
rect 13570 39919 13586 39983
rect 13650 39919 13666 39983
rect 13730 39919 13746 39983
rect 13810 39919 13826 39983
rect 13890 39919 13906 39983
rect 13970 39919 13986 39983
rect 14050 39919 14066 39983
rect 14130 39919 14146 39983
rect 14210 39919 14226 39983
rect 14290 39919 14306 39983
rect 14370 39919 14386 39983
rect 14450 39919 14466 39983
rect 14530 39919 14546 39983
rect 14610 39919 14626 39983
rect 14690 39919 14706 39983
rect 14770 39919 14786 39983
rect 14850 39919 14858 39983
rect 12264 39902 14858 39919
rect 12264 39838 12306 39902
rect 12370 39838 12386 39902
rect 12450 39838 12466 39902
rect 12530 39838 12546 39902
rect 12610 39838 12626 39902
rect 12690 39838 12706 39902
rect 12770 39838 12786 39902
rect 12850 39838 12866 39902
rect 12930 39838 12946 39902
rect 13010 39838 13026 39902
rect 13090 39838 13106 39902
rect 13170 39838 13186 39902
rect 13250 39838 13266 39902
rect 13330 39838 13346 39902
rect 13410 39838 13426 39902
rect 13490 39838 13506 39902
rect 13570 39838 13586 39902
rect 13650 39838 13666 39902
rect 13730 39838 13746 39902
rect 13810 39838 13826 39902
rect 13890 39838 13906 39902
rect 13970 39838 13986 39902
rect 14050 39838 14066 39902
rect 14130 39838 14146 39902
rect 14210 39838 14226 39902
rect 14290 39838 14306 39902
rect 14370 39838 14386 39902
rect 14450 39838 14466 39902
rect 14530 39838 14546 39902
rect 14610 39838 14626 39902
rect 14690 39838 14706 39902
rect 14770 39838 14786 39902
rect 14850 39838 14858 39902
rect 12264 39821 14858 39838
rect 12264 39757 12306 39821
rect 12370 39757 12386 39821
rect 12450 39757 12466 39821
rect 12530 39757 12546 39821
rect 12610 39757 12626 39821
rect 12690 39757 12706 39821
rect 12770 39757 12786 39821
rect 12850 39757 12866 39821
rect 12930 39757 12946 39821
rect 13010 39757 13026 39821
rect 13090 39757 13106 39821
rect 13170 39757 13186 39821
rect 13250 39757 13266 39821
rect 13330 39757 13346 39821
rect 13410 39757 13426 39821
rect 13490 39757 13506 39821
rect 13570 39757 13586 39821
rect 13650 39757 13666 39821
rect 13730 39757 13746 39821
rect 13810 39757 13826 39821
rect 13890 39757 13906 39821
rect 13970 39757 13986 39821
rect 14050 39757 14066 39821
rect 14130 39757 14146 39821
rect 14210 39757 14226 39821
rect 14290 39757 14306 39821
rect 14370 39757 14386 39821
rect 14450 39757 14466 39821
rect 14530 39757 14546 39821
rect 14610 39757 14626 39821
rect 14690 39757 14706 39821
rect 14770 39757 14786 39821
rect 14850 39757 14858 39821
rect 12264 39740 14858 39757
rect 12264 39676 12306 39740
rect 12370 39676 12386 39740
rect 12450 39676 12466 39740
rect 12530 39676 12546 39740
rect 12610 39676 12626 39740
rect 12690 39676 12706 39740
rect 12770 39676 12786 39740
rect 12850 39676 12866 39740
rect 12930 39676 12946 39740
rect 13010 39676 13026 39740
rect 13090 39676 13106 39740
rect 13170 39676 13186 39740
rect 13250 39676 13266 39740
rect 13330 39676 13346 39740
rect 13410 39676 13426 39740
rect 13490 39676 13506 39740
rect 13570 39676 13586 39740
rect 13650 39676 13666 39740
rect 13730 39676 13746 39740
rect 13810 39676 13826 39740
rect 13890 39676 13906 39740
rect 13970 39676 13986 39740
rect 14050 39676 14066 39740
rect 14130 39676 14146 39740
rect 14210 39676 14226 39740
rect 14290 39676 14306 39740
rect 14370 39676 14386 39740
rect 14450 39676 14466 39740
rect 14530 39676 14546 39740
rect 14610 39676 14626 39740
rect 14690 39676 14706 39740
rect 14770 39676 14786 39740
rect 14850 39676 14858 39740
rect 12264 39659 14858 39676
rect 12264 39595 12306 39659
rect 12370 39595 12386 39659
rect 12450 39595 12466 39659
rect 12530 39595 12546 39659
rect 12610 39595 12626 39659
rect 12690 39595 12706 39659
rect 12770 39595 12786 39659
rect 12850 39595 12866 39659
rect 12930 39595 12946 39659
rect 13010 39595 13026 39659
rect 13090 39595 13106 39659
rect 13170 39595 13186 39659
rect 13250 39595 13266 39659
rect 13330 39595 13346 39659
rect 13410 39595 13426 39659
rect 13490 39595 13506 39659
rect 13570 39595 13586 39659
rect 13650 39595 13666 39659
rect 13730 39595 13746 39659
rect 13810 39595 13826 39659
rect 13890 39595 13906 39659
rect 13970 39595 13986 39659
rect 14050 39595 14066 39659
rect 14130 39595 14146 39659
rect 14210 39595 14226 39659
rect 14290 39595 14306 39659
rect 14370 39595 14386 39659
rect 14450 39595 14466 39659
rect 14530 39595 14546 39659
rect 14610 39595 14626 39659
rect 14690 39595 14706 39659
rect 14770 39595 14786 39659
rect 14850 39595 14858 39659
rect 12264 39578 14858 39595
rect 12264 39514 12306 39578
rect 12370 39514 12386 39578
rect 12450 39514 12466 39578
rect 12530 39514 12546 39578
rect 12610 39514 12626 39578
rect 12690 39514 12706 39578
rect 12770 39514 12786 39578
rect 12850 39514 12866 39578
rect 12930 39514 12946 39578
rect 13010 39514 13026 39578
rect 13090 39514 13106 39578
rect 13170 39514 13186 39578
rect 13250 39514 13266 39578
rect 13330 39514 13346 39578
rect 13410 39514 13426 39578
rect 13490 39514 13506 39578
rect 13570 39514 13586 39578
rect 13650 39514 13666 39578
rect 13730 39514 13746 39578
rect 13810 39514 13826 39578
rect 13890 39514 13906 39578
rect 13970 39514 13986 39578
rect 14050 39514 14066 39578
rect 14130 39514 14146 39578
rect 14210 39514 14226 39578
rect 14290 39514 14306 39578
rect 14370 39514 14386 39578
rect 14450 39514 14466 39578
rect 14530 39514 14546 39578
rect 14610 39514 14626 39578
rect 14690 39514 14706 39578
rect 14770 39514 14786 39578
rect 14850 39514 14858 39578
rect 12264 39497 14858 39514
rect 12264 39438 12306 39497
rect 2669 39435 12306 39438
rect 2669 39433 3031 39435
rect 99 39416 3031 39433
rect 99 39352 125 39416
rect 189 39352 205 39416
rect 269 39352 285 39416
rect 349 39352 365 39416
rect 429 39352 445 39416
rect 509 39352 525 39416
rect 589 39352 605 39416
rect 669 39352 685 39416
rect 749 39352 765 39416
rect 829 39352 845 39416
rect 909 39352 925 39416
rect 989 39352 1005 39416
rect 1069 39352 1085 39416
rect 1149 39352 1165 39416
rect 1229 39352 1245 39416
rect 1309 39352 1325 39416
rect 1389 39352 1405 39416
rect 1469 39352 1485 39416
rect 1549 39352 1565 39416
rect 1629 39352 1645 39416
rect 1709 39352 1725 39416
rect 1789 39352 1805 39416
rect 1869 39352 1885 39416
rect 1949 39352 1965 39416
rect 2029 39352 2045 39416
rect 2109 39352 2125 39416
rect 2189 39352 2205 39416
rect 2269 39352 2285 39416
rect 2349 39352 2365 39416
rect 2429 39352 2445 39416
rect 2509 39352 2525 39416
rect 2589 39352 2605 39416
rect 2669 39399 3031 39416
tri 3031 39399 3067 39435 nw
tri 11927 39399 11963 39435 ne
rect 11963 39433 12306 39435
rect 12370 39433 12386 39497
rect 12450 39433 12466 39497
rect 12530 39433 12546 39497
rect 12610 39433 12626 39497
rect 12690 39433 12706 39497
rect 12770 39433 12786 39497
rect 12850 39433 12866 39497
rect 12930 39433 12946 39497
rect 13010 39433 13026 39497
rect 13090 39433 13106 39497
rect 13170 39433 13186 39497
rect 13250 39433 13266 39497
rect 13330 39433 13346 39497
rect 13410 39433 13426 39497
rect 13490 39433 13506 39497
rect 13570 39433 13586 39497
rect 13650 39433 13666 39497
rect 13730 39433 13746 39497
rect 13810 39433 13826 39497
rect 13890 39433 13906 39497
rect 13970 39433 13986 39497
rect 14050 39433 14066 39497
rect 14130 39433 14146 39497
rect 14210 39433 14226 39497
rect 14290 39433 14306 39497
rect 14370 39433 14386 39497
rect 14450 39433 14466 39497
rect 14530 39433 14546 39497
rect 14610 39433 14626 39497
rect 14690 39433 14706 39497
rect 14770 39433 14786 39497
rect 14850 39433 14858 39497
rect 11963 39416 14858 39433
rect 11963 39399 12306 39416
rect 2669 39393 2873 39399
rect 2669 39352 2753 39393
rect 99 39335 2753 39352
rect 99 39271 125 39335
rect 189 39271 205 39335
rect 269 39271 285 39335
rect 349 39271 365 39335
rect 429 39271 445 39335
rect 509 39271 525 39335
rect 589 39271 605 39335
rect 669 39271 685 39335
rect 749 39271 765 39335
rect 829 39271 845 39335
rect 909 39271 925 39335
rect 989 39271 1005 39335
rect 1069 39271 1085 39335
rect 1149 39271 1165 39335
rect 1229 39271 1245 39335
rect 1309 39271 1325 39335
rect 1389 39271 1405 39335
rect 1469 39271 1485 39335
rect 1549 39271 1565 39335
rect 1629 39271 1645 39335
rect 1709 39271 1725 39335
rect 1789 39271 1805 39335
rect 1869 39271 1885 39335
rect 1949 39271 1965 39335
rect 2029 39271 2045 39335
rect 2109 39271 2125 39335
rect 2189 39271 2205 39335
rect 2269 39271 2285 39335
rect 2349 39271 2365 39335
rect 2429 39271 2445 39335
rect 2509 39271 2525 39335
rect 2589 39271 2605 39335
rect 2669 39329 2753 39335
rect 2817 39329 2873 39393
rect 2669 39311 2873 39329
rect 2669 39271 2753 39311
rect 99 39254 2753 39271
rect 99 39190 125 39254
rect 189 39190 205 39254
rect 269 39190 285 39254
rect 349 39190 365 39254
rect 429 39190 445 39254
rect 509 39190 525 39254
rect 589 39190 605 39254
rect 669 39190 685 39254
rect 749 39190 765 39254
rect 829 39190 845 39254
rect 909 39190 925 39254
rect 989 39190 1005 39254
rect 1069 39190 1085 39254
rect 1149 39190 1165 39254
rect 1229 39190 1245 39254
rect 1309 39190 1325 39254
rect 1389 39190 1405 39254
rect 1469 39190 1485 39254
rect 1549 39190 1565 39254
rect 1629 39190 1645 39254
rect 1709 39190 1725 39254
rect 1789 39190 1805 39254
rect 1869 39190 1885 39254
rect 1949 39190 1965 39254
rect 2029 39190 2045 39254
rect 2109 39190 2125 39254
rect 2189 39190 2205 39254
rect 2269 39190 2285 39254
rect 2349 39190 2365 39254
rect 2429 39190 2445 39254
rect 2509 39190 2525 39254
rect 2589 39190 2605 39254
rect 2669 39247 2753 39254
rect 2817 39247 2873 39311
rect 2669 39241 2873 39247
tri 2873 39241 3031 39399 nw
tri 11963 39241 12121 39399 ne
rect 12121 39393 12306 39399
rect 12121 39329 12170 39393
rect 12234 39352 12306 39393
rect 12370 39352 12386 39416
rect 12450 39352 12466 39416
rect 12530 39352 12546 39416
rect 12610 39352 12626 39416
rect 12690 39352 12706 39416
rect 12770 39352 12786 39416
rect 12850 39352 12866 39416
rect 12930 39352 12946 39416
rect 13010 39352 13026 39416
rect 13090 39352 13106 39416
rect 13170 39352 13186 39416
rect 13250 39352 13266 39416
rect 13330 39352 13346 39416
rect 13410 39352 13426 39416
rect 13490 39352 13506 39416
rect 13570 39352 13586 39416
rect 13650 39352 13666 39416
rect 13730 39352 13746 39416
rect 13810 39352 13826 39416
rect 13890 39352 13906 39416
rect 13970 39352 13986 39416
rect 14050 39352 14066 39416
rect 14130 39352 14146 39416
rect 14210 39352 14226 39416
rect 14290 39352 14306 39416
rect 14370 39352 14386 39416
rect 14450 39352 14466 39416
rect 14530 39352 14546 39416
rect 14610 39352 14626 39416
rect 14690 39352 14706 39416
rect 14770 39352 14786 39416
rect 14850 39352 14858 39416
rect 12234 39335 14858 39352
rect 12234 39329 12306 39335
rect 12121 39311 12306 39329
rect 12121 39247 12170 39311
rect 12234 39271 12306 39311
rect 12370 39271 12386 39335
rect 12450 39271 12466 39335
rect 12530 39271 12546 39335
rect 12610 39271 12626 39335
rect 12690 39271 12706 39335
rect 12770 39271 12786 39335
rect 12850 39271 12866 39335
rect 12930 39271 12946 39335
rect 13010 39271 13026 39335
rect 13090 39271 13106 39335
rect 13170 39271 13186 39335
rect 13250 39271 13266 39335
rect 13330 39271 13346 39335
rect 13410 39271 13426 39335
rect 13490 39271 13506 39335
rect 13570 39271 13586 39335
rect 13650 39271 13666 39335
rect 13730 39271 13746 39335
rect 13810 39271 13826 39335
rect 13890 39271 13906 39335
rect 13970 39271 13986 39335
rect 14050 39271 14066 39335
rect 14130 39271 14146 39335
rect 14210 39271 14226 39335
rect 14290 39271 14306 39335
rect 14370 39271 14386 39335
rect 14450 39271 14466 39335
rect 14530 39271 14546 39335
rect 14610 39271 14626 39335
rect 14690 39271 14706 39335
rect 14770 39271 14786 39335
rect 14850 39271 14858 39335
rect 12234 39254 14858 39271
rect 12234 39247 12306 39254
rect 12121 39241 12306 39247
rect 2669 39190 2700 39241
rect 99 39173 2700 39190
rect 99 39109 125 39173
rect 189 39109 205 39173
rect 269 39109 285 39173
rect 349 39109 365 39173
rect 429 39109 445 39173
rect 509 39109 525 39173
rect 589 39109 605 39173
rect 669 39109 685 39173
rect 749 39109 765 39173
rect 829 39109 845 39173
rect 909 39109 925 39173
rect 989 39109 1005 39173
rect 1069 39109 1085 39173
rect 1149 39109 1165 39173
rect 1229 39109 1245 39173
rect 1309 39109 1325 39173
rect 1389 39109 1405 39173
rect 1469 39109 1485 39173
rect 1549 39109 1565 39173
rect 1629 39109 1645 39173
rect 1709 39109 1725 39173
rect 1789 39109 1805 39173
rect 1869 39109 1885 39173
rect 1949 39109 1965 39173
rect 2029 39109 2045 39173
rect 2109 39109 2125 39173
rect 2189 39109 2205 39173
rect 2269 39109 2285 39173
rect 2349 39109 2365 39173
rect 2429 39109 2445 39173
rect 2509 39109 2525 39173
rect 2589 39109 2605 39173
rect 2669 39109 2700 39173
rect 99 39092 2700 39109
rect 99 39028 125 39092
rect 189 39028 205 39092
rect 269 39028 285 39092
rect 349 39028 365 39092
rect 429 39028 445 39092
rect 509 39028 525 39092
rect 589 39028 605 39092
rect 669 39028 685 39092
rect 749 39028 765 39092
rect 829 39028 845 39092
rect 909 39028 925 39092
rect 989 39028 1005 39092
rect 1069 39028 1085 39092
rect 1149 39028 1165 39092
rect 1229 39028 1245 39092
rect 1309 39028 1325 39092
rect 1389 39028 1405 39092
rect 1469 39028 1485 39092
rect 1549 39028 1565 39092
rect 1629 39028 1645 39092
rect 1709 39028 1725 39092
rect 1789 39028 1805 39092
rect 1869 39028 1885 39092
rect 1949 39028 1965 39092
rect 2029 39028 2045 39092
rect 2109 39028 2125 39092
rect 2189 39028 2205 39092
rect 2269 39028 2285 39092
rect 2349 39028 2365 39092
rect 2429 39028 2445 39092
rect 2509 39028 2525 39092
rect 2589 39028 2605 39092
rect 2669 39028 2700 39092
tri 2700 39068 2873 39241 nw
tri 12121 39068 12294 39241 ne
rect 12294 39190 12306 39241
rect 12370 39190 12386 39254
rect 12450 39190 12466 39254
rect 12530 39190 12546 39254
rect 12610 39190 12626 39254
rect 12690 39190 12706 39254
rect 12770 39190 12786 39254
rect 12850 39190 12866 39254
rect 12930 39190 12946 39254
rect 13010 39190 13026 39254
rect 13090 39190 13106 39254
rect 13170 39190 13186 39254
rect 13250 39190 13266 39254
rect 13330 39190 13346 39254
rect 13410 39190 13426 39254
rect 13490 39190 13506 39254
rect 13570 39190 13586 39254
rect 13650 39190 13666 39254
rect 13730 39190 13746 39254
rect 13810 39190 13826 39254
rect 13890 39190 13906 39254
rect 13970 39190 13986 39254
rect 14050 39190 14066 39254
rect 14130 39190 14146 39254
rect 14210 39190 14226 39254
rect 14290 39190 14306 39254
rect 14370 39190 14386 39254
rect 14450 39190 14466 39254
rect 14530 39190 14546 39254
rect 14610 39190 14626 39254
rect 14690 39190 14706 39254
rect 14770 39190 14786 39254
rect 14850 39190 14858 39254
rect 12294 39173 14858 39190
rect 12294 39109 12306 39173
rect 12370 39109 12386 39173
rect 12450 39109 12466 39173
rect 12530 39109 12546 39173
rect 12610 39109 12626 39173
rect 12690 39109 12706 39173
rect 12770 39109 12786 39173
rect 12850 39109 12866 39173
rect 12930 39109 12946 39173
rect 13010 39109 13026 39173
rect 13090 39109 13106 39173
rect 13170 39109 13186 39173
rect 13250 39109 13266 39173
rect 13330 39109 13346 39173
rect 13410 39109 13426 39173
rect 13490 39109 13506 39173
rect 13570 39109 13586 39173
rect 13650 39109 13666 39173
rect 13730 39109 13746 39173
rect 13810 39109 13826 39173
rect 13890 39109 13906 39173
rect 13970 39109 13986 39173
rect 14050 39109 14066 39173
rect 14130 39109 14146 39173
rect 14210 39109 14226 39173
rect 14290 39109 14306 39173
rect 14370 39109 14386 39173
rect 14450 39109 14466 39173
rect 14530 39109 14546 39173
rect 14610 39109 14626 39173
rect 14690 39109 14706 39173
rect 14770 39109 14786 39173
rect 14850 39109 14858 39173
rect 12294 39092 14858 39109
rect 12294 39068 12306 39092
tri 12294 39062 12300 39068 ne
rect 99 39011 2700 39028
rect 99 35187 125 39011
rect 2669 35187 2700 39011
rect 99 34631 2700 35187
rect 12300 39028 12306 39068
rect 12370 39028 12386 39092
rect 12450 39028 12466 39092
rect 12530 39028 12546 39092
rect 12610 39028 12626 39092
rect 12690 39028 12706 39092
rect 12770 39028 12786 39092
rect 12850 39028 12866 39092
rect 12930 39028 12946 39092
rect 13010 39028 13026 39092
rect 13090 39028 13106 39092
rect 13170 39028 13186 39092
rect 13250 39028 13266 39092
rect 13330 39028 13346 39092
rect 13410 39028 13426 39092
rect 13490 39028 13506 39092
rect 13570 39028 13586 39092
rect 13650 39028 13666 39092
rect 13730 39028 13746 39092
rect 13810 39028 13826 39092
rect 13890 39028 13906 39092
rect 13970 39028 13986 39092
rect 14050 39028 14066 39092
rect 14130 39028 14146 39092
rect 14210 39028 14226 39092
rect 14290 39028 14306 39092
rect 14370 39028 14386 39092
rect 14450 39028 14466 39092
rect 14530 39028 14546 39092
rect 14610 39028 14626 39092
rect 14690 39028 14706 39092
rect 14770 39028 14786 39092
rect 14850 39028 14858 39092
rect 12300 39011 14858 39028
rect 12300 35187 12306 39011
rect 14850 35187 14858 39011
rect 12300 34664 14858 35187
rect 104 12534 4874 12536
rect 104 12470 105 12534
rect 169 12470 187 12534
rect 251 12470 269 12534
rect 333 12470 351 12534
rect 415 12470 433 12534
rect 497 12470 515 12534
rect 579 12470 597 12534
rect 661 12470 678 12534
rect 742 12470 759 12534
rect 823 12470 840 12534
rect 904 12470 921 12534
rect 985 12470 1002 12534
rect 1066 12470 1083 12534
rect 1147 12470 1164 12534
rect 1228 12470 1245 12534
rect 1309 12470 1326 12534
rect 1390 12470 1407 12534
rect 1471 12470 1488 12534
rect 1552 12470 1569 12534
rect 1633 12470 1650 12534
rect 1714 12470 1731 12534
rect 1795 12470 1812 12534
rect 1876 12470 1893 12534
rect 1957 12470 1974 12534
rect 2038 12470 2055 12534
rect 2119 12470 2136 12534
rect 2200 12470 2217 12534
rect 2281 12470 2298 12534
rect 2362 12470 2379 12534
rect 2443 12470 2460 12534
rect 2524 12470 2541 12534
rect 2605 12470 2622 12534
rect 2686 12470 2703 12534
rect 2767 12470 2784 12534
rect 2848 12470 2865 12534
rect 2929 12470 2946 12534
rect 3010 12470 3027 12534
rect 3091 12470 3108 12534
rect 3172 12470 3189 12534
rect 3253 12470 3270 12534
rect 3334 12470 3351 12534
rect 3415 12470 3432 12534
rect 3496 12470 3513 12534
rect 3577 12470 3594 12534
rect 3658 12470 3675 12534
rect 3739 12470 3756 12534
rect 3820 12470 3837 12534
rect 3901 12470 3918 12534
rect 3982 12470 3999 12534
rect 4063 12470 4080 12534
rect 4144 12470 4161 12534
rect 4225 12470 4242 12534
rect 4306 12470 4323 12534
rect 4387 12470 4404 12534
rect 4468 12470 4485 12534
rect 4549 12470 4566 12534
rect 4630 12470 4647 12534
rect 4711 12470 4728 12534
rect 4792 12470 4809 12534
rect 4873 12470 4874 12534
rect 104 12452 4874 12470
rect 104 12388 105 12452
rect 169 12388 187 12452
rect 251 12388 269 12452
rect 333 12388 351 12452
rect 415 12388 433 12452
rect 497 12388 515 12452
rect 579 12388 597 12452
rect 661 12388 678 12452
rect 742 12388 759 12452
rect 823 12388 840 12452
rect 904 12388 921 12452
rect 985 12388 1002 12452
rect 1066 12388 1083 12452
rect 1147 12388 1164 12452
rect 1228 12388 1245 12452
rect 1309 12388 1326 12452
rect 1390 12388 1407 12452
rect 1471 12388 1488 12452
rect 1552 12388 1569 12452
rect 1633 12388 1650 12452
rect 1714 12388 1731 12452
rect 1795 12388 1812 12452
rect 1876 12388 1893 12452
rect 1957 12388 1974 12452
rect 2038 12388 2055 12452
rect 2119 12388 2136 12452
rect 2200 12388 2217 12452
rect 2281 12388 2298 12452
rect 2362 12388 2379 12452
rect 2443 12388 2460 12452
rect 2524 12388 2541 12452
rect 2605 12388 2622 12452
rect 2686 12388 2703 12452
rect 2767 12388 2784 12452
rect 2848 12388 2865 12452
rect 2929 12388 2946 12452
rect 3010 12388 3027 12452
rect 3091 12388 3108 12452
rect 3172 12388 3189 12452
rect 3253 12388 3270 12452
rect 3334 12388 3351 12452
rect 3415 12388 3432 12452
rect 3496 12388 3513 12452
rect 3577 12388 3594 12452
rect 3658 12388 3675 12452
rect 3739 12388 3756 12452
rect 3820 12388 3837 12452
rect 3901 12388 3918 12452
rect 3982 12388 3999 12452
rect 4063 12388 4080 12452
rect 4144 12388 4161 12452
rect 4225 12388 4242 12452
rect 4306 12388 4323 12452
rect 4387 12388 4404 12452
rect 4468 12388 4485 12452
rect 4549 12388 4566 12452
rect 4630 12388 4647 12452
rect 4711 12388 4728 12452
rect 4792 12388 4809 12452
rect 4873 12388 4874 12452
rect 104 12370 4874 12388
rect 104 12306 105 12370
rect 169 12306 187 12370
rect 251 12306 269 12370
rect 333 12306 351 12370
rect 415 12306 433 12370
rect 497 12306 515 12370
rect 579 12306 597 12370
rect 661 12306 678 12370
rect 742 12306 759 12370
rect 823 12306 840 12370
rect 904 12306 921 12370
rect 985 12306 1002 12370
rect 1066 12306 1083 12370
rect 1147 12306 1164 12370
rect 1228 12306 1245 12370
rect 1309 12306 1326 12370
rect 1390 12306 1407 12370
rect 1471 12306 1488 12370
rect 1552 12306 1569 12370
rect 1633 12306 1650 12370
rect 1714 12306 1731 12370
rect 1795 12306 1812 12370
rect 1876 12306 1893 12370
rect 1957 12306 1974 12370
rect 2038 12306 2055 12370
rect 2119 12306 2136 12370
rect 2200 12306 2217 12370
rect 2281 12306 2298 12370
rect 2362 12306 2379 12370
rect 2443 12306 2460 12370
rect 2524 12306 2541 12370
rect 2605 12306 2622 12370
rect 2686 12306 2703 12370
rect 2767 12306 2784 12370
rect 2848 12306 2865 12370
rect 2929 12306 2946 12370
rect 3010 12306 3027 12370
rect 3091 12306 3108 12370
rect 3172 12306 3189 12370
rect 3253 12306 3270 12370
rect 3334 12306 3351 12370
rect 3415 12306 3432 12370
rect 3496 12306 3513 12370
rect 3577 12306 3594 12370
rect 3658 12306 3675 12370
rect 3739 12306 3756 12370
rect 3820 12306 3837 12370
rect 3901 12306 3918 12370
rect 3982 12306 3999 12370
rect 4063 12306 4080 12370
rect 4144 12306 4161 12370
rect 4225 12306 4242 12370
rect 4306 12306 4323 12370
rect 4387 12306 4404 12370
rect 4468 12306 4485 12370
rect 4549 12306 4566 12370
rect 4630 12306 4647 12370
rect 4711 12306 4728 12370
rect 4792 12306 4809 12370
rect 4873 12306 4874 12370
rect 104 12288 4874 12306
rect 104 12224 105 12288
rect 169 12224 187 12288
rect 251 12224 269 12288
rect 333 12224 351 12288
rect 415 12224 433 12288
rect 497 12224 515 12288
rect 579 12224 597 12288
rect 661 12224 678 12288
rect 742 12224 759 12288
rect 823 12224 840 12288
rect 904 12224 921 12288
rect 985 12224 1002 12288
rect 1066 12224 1083 12288
rect 1147 12224 1164 12288
rect 1228 12224 1245 12288
rect 1309 12224 1326 12288
rect 1390 12224 1407 12288
rect 1471 12224 1488 12288
rect 1552 12224 1569 12288
rect 1633 12224 1650 12288
rect 1714 12224 1731 12288
rect 1795 12224 1812 12288
rect 1876 12224 1893 12288
rect 1957 12224 1974 12288
rect 2038 12224 2055 12288
rect 2119 12224 2136 12288
rect 2200 12224 2217 12288
rect 2281 12224 2298 12288
rect 2362 12224 2379 12288
rect 2443 12224 2460 12288
rect 2524 12224 2541 12288
rect 2605 12224 2622 12288
rect 2686 12224 2703 12288
rect 2767 12224 2784 12288
rect 2848 12224 2865 12288
rect 2929 12224 2946 12288
rect 3010 12224 3027 12288
rect 3091 12224 3108 12288
rect 3172 12224 3189 12288
rect 3253 12224 3270 12288
rect 3334 12224 3351 12288
rect 3415 12224 3432 12288
rect 3496 12224 3513 12288
rect 3577 12224 3594 12288
rect 3658 12224 3675 12288
rect 3739 12224 3756 12288
rect 3820 12224 3837 12288
rect 3901 12224 3918 12288
rect 3982 12224 3999 12288
rect 4063 12224 4080 12288
rect 4144 12224 4161 12288
rect 4225 12224 4242 12288
rect 4306 12224 4323 12288
rect 4387 12224 4404 12288
rect 4468 12224 4485 12288
rect 4549 12224 4566 12288
rect 4630 12224 4647 12288
rect 4711 12224 4728 12288
rect 4792 12224 4809 12288
rect 4873 12224 4874 12288
rect 104 12206 4874 12224
rect 104 12142 105 12206
rect 169 12142 187 12206
rect 251 12142 269 12206
rect 333 12142 351 12206
rect 415 12142 433 12206
rect 497 12142 515 12206
rect 579 12142 597 12206
rect 661 12142 678 12206
rect 742 12142 759 12206
rect 823 12142 840 12206
rect 904 12142 921 12206
rect 985 12142 1002 12206
rect 1066 12142 1083 12206
rect 1147 12142 1164 12206
rect 1228 12142 1245 12206
rect 1309 12142 1326 12206
rect 1390 12142 1407 12206
rect 1471 12142 1488 12206
rect 1552 12142 1569 12206
rect 1633 12142 1650 12206
rect 1714 12142 1731 12206
rect 1795 12142 1812 12206
rect 1876 12142 1893 12206
rect 1957 12142 1974 12206
rect 2038 12142 2055 12206
rect 2119 12142 2136 12206
rect 2200 12142 2217 12206
rect 2281 12142 2298 12206
rect 2362 12142 2379 12206
rect 2443 12142 2460 12206
rect 2524 12142 2541 12206
rect 2605 12142 2622 12206
rect 2686 12142 2703 12206
rect 2767 12142 2784 12206
rect 2848 12142 2865 12206
rect 2929 12142 2946 12206
rect 3010 12142 3027 12206
rect 3091 12142 3108 12206
rect 3172 12142 3189 12206
rect 3253 12142 3270 12206
rect 3334 12142 3351 12206
rect 3415 12142 3432 12206
rect 3496 12142 3513 12206
rect 3577 12142 3594 12206
rect 3658 12142 3675 12206
rect 3739 12142 3756 12206
rect 3820 12142 3837 12206
rect 3901 12142 3918 12206
rect 3982 12142 3999 12206
rect 4063 12142 4080 12206
rect 4144 12142 4161 12206
rect 4225 12142 4242 12206
rect 4306 12142 4323 12206
rect 4387 12142 4404 12206
rect 4468 12142 4485 12206
rect 4549 12142 4566 12206
rect 4630 12142 4647 12206
rect 4711 12142 4728 12206
rect 4792 12142 4809 12206
rect 4873 12142 4874 12206
rect 104 12124 4874 12142
rect 104 12060 105 12124
rect 169 12060 187 12124
rect 251 12060 269 12124
rect 333 12060 351 12124
rect 415 12060 433 12124
rect 497 12060 515 12124
rect 579 12060 597 12124
rect 661 12060 678 12124
rect 742 12060 759 12124
rect 823 12060 840 12124
rect 904 12060 921 12124
rect 985 12060 1002 12124
rect 1066 12060 1083 12124
rect 1147 12060 1164 12124
rect 1228 12060 1245 12124
rect 1309 12060 1326 12124
rect 1390 12060 1407 12124
rect 1471 12060 1488 12124
rect 1552 12060 1569 12124
rect 1633 12060 1650 12124
rect 1714 12060 1731 12124
rect 1795 12060 1812 12124
rect 1876 12060 1893 12124
rect 1957 12060 1974 12124
rect 2038 12060 2055 12124
rect 2119 12060 2136 12124
rect 2200 12060 2217 12124
rect 2281 12060 2298 12124
rect 2362 12060 2379 12124
rect 2443 12060 2460 12124
rect 2524 12060 2541 12124
rect 2605 12060 2622 12124
rect 2686 12060 2703 12124
rect 2767 12060 2784 12124
rect 2848 12060 2865 12124
rect 2929 12060 2946 12124
rect 3010 12060 3027 12124
rect 3091 12060 3108 12124
rect 3172 12060 3189 12124
rect 3253 12060 3270 12124
rect 3334 12060 3351 12124
rect 3415 12060 3432 12124
rect 3496 12060 3513 12124
rect 3577 12060 3594 12124
rect 3658 12060 3675 12124
rect 3739 12060 3756 12124
rect 3820 12060 3837 12124
rect 3901 12060 3918 12124
rect 3982 12060 3999 12124
rect 4063 12060 4080 12124
rect 4144 12060 4161 12124
rect 4225 12060 4242 12124
rect 4306 12060 4323 12124
rect 4387 12060 4404 12124
rect 4468 12060 4485 12124
rect 4549 12060 4566 12124
rect 4630 12060 4647 12124
rect 4711 12060 4728 12124
rect 4792 12060 4809 12124
rect 4873 12060 4874 12124
rect 104 12042 4874 12060
rect 104 11978 105 12042
rect 169 11978 187 12042
rect 251 11978 269 12042
rect 333 11978 351 12042
rect 415 11978 433 12042
rect 497 11978 515 12042
rect 579 11978 597 12042
rect 661 11978 678 12042
rect 742 11978 759 12042
rect 823 11978 840 12042
rect 904 11978 921 12042
rect 985 11978 1002 12042
rect 1066 11978 1083 12042
rect 1147 11978 1164 12042
rect 1228 11978 1245 12042
rect 1309 11978 1326 12042
rect 1390 11978 1407 12042
rect 1471 11978 1488 12042
rect 1552 11978 1569 12042
rect 1633 11978 1650 12042
rect 1714 11978 1731 12042
rect 1795 11978 1812 12042
rect 1876 11978 1893 12042
rect 1957 11978 1974 12042
rect 2038 11978 2055 12042
rect 2119 11978 2136 12042
rect 2200 11978 2217 12042
rect 2281 11978 2298 12042
rect 2362 11978 2379 12042
rect 2443 11978 2460 12042
rect 2524 11978 2541 12042
rect 2605 11978 2622 12042
rect 2686 11978 2703 12042
rect 2767 11978 2784 12042
rect 2848 11978 2865 12042
rect 2929 11978 2946 12042
rect 3010 11978 3027 12042
rect 3091 11978 3108 12042
rect 3172 11978 3189 12042
rect 3253 11978 3270 12042
rect 3334 11978 3351 12042
rect 3415 11978 3432 12042
rect 3496 11978 3513 12042
rect 3577 11978 3594 12042
rect 3658 11978 3675 12042
rect 3739 11978 3756 12042
rect 3820 11978 3837 12042
rect 3901 11978 3918 12042
rect 3982 11978 3999 12042
rect 4063 11978 4080 12042
rect 4144 11978 4161 12042
rect 4225 11978 4242 12042
rect 4306 11978 4323 12042
rect 4387 11978 4404 12042
rect 4468 11978 4485 12042
rect 4549 11978 4566 12042
rect 4630 11978 4647 12042
rect 4711 11978 4728 12042
rect 4792 11978 4809 12042
rect 4873 11978 4874 12042
rect 104 11960 4874 11978
rect 104 11896 105 11960
rect 169 11896 187 11960
rect 251 11896 269 11960
rect 333 11896 351 11960
rect 415 11896 433 11960
rect 497 11896 515 11960
rect 579 11896 597 11960
rect 661 11896 678 11960
rect 742 11896 759 11960
rect 823 11896 840 11960
rect 904 11896 921 11960
rect 985 11896 1002 11960
rect 1066 11896 1083 11960
rect 1147 11896 1164 11960
rect 1228 11896 1245 11960
rect 1309 11896 1326 11960
rect 1390 11896 1407 11960
rect 1471 11896 1488 11960
rect 1552 11896 1569 11960
rect 1633 11896 1650 11960
rect 1714 11896 1731 11960
rect 1795 11896 1812 11960
rect 1876 11896 1893 11960
rect 1957 11896 1974 11960
rect 2038 11896 2055 11960
rect 2119 11896 2136 11960
rect 2200 11896 2217 11960
rect 2281 11896 2298 11960
rect 2362 11896 2379 11960
rect 2443 11896 2460 11960
rect 2524 11896 2541 11960
rect 2605 11896 2622 11960
rect 2686 11896 2703 11960
rect 2767 11896 2784 11960
rect 2848 11896 2865 11960
rect 2929 11896 2946 11960
rect 3010 11896 3027 11960
rect 3091 11896 3108 11960
rect 3172 11896 3189 11960
rect 3253 11896 3270 11960
rect 3334 11896 3351 11960
rect 3415 11896 3432 11960
rect 3496 11896 3513 11960
rect 3577 11896 3594 11960
rect 3658 11896 3675 11960
rect 3739 11896 3756 11960
rect 3820 11896 3837 11960
rect 3901 11896 3918 11960
rect 3982 11896 3999 11960
rect 4063 11896 4080 11960
rect 4144 11896 4161 11960
rect 4225 11896 4242 11960
rect 4306 11896 4323 11960
rect 4387 11896 4404 11960
rect 4468 11896 4485 11960
rect 4549 11896 4566 11960
rect 4630 11896 4647 11960
rect 4711 11896 4728 11960
rect 4792 11896 4809 11960
rect 4873 11896 4874 11960
rect 104 11878 4874 11896
rect 104 11814 105 11878
rect 169 11814 187 11878
rect 251 11814 269 11878
rect 333 11814 351 11878
rect 415 11814 433 11878
rect 497 11814 515 11878
rect 579 11814 597 11878
rect 661 11814 678 11878
rect 742 11814 759 11878
rect 823 11814 840 11878
rect 904 11814 921 11878
rect 985 11814 1002 11878
rect 1066 11814 1083 11878
rect 1147 11814 1164 11878
rect 1228 11814 1245 11878
rect 1309 11814 1326 11878
rect 1390 11814 1407 11878
rect 1471 11814 1488 11878
rect 1552 11814 1569 11878
rect 1633 11814 1650 11878
rect 1714 11814 1731 11878
rect 1795 11814 1812 11878
rect 1876 11814 1893 11878
rect 1957 11814 1974 11878
rect 2038 11814 2055 11878
rect 2119 11814 2136 11878
rect 2200 11814 2217 11878
rect 2281 11814 2298 11878
rect 2362 11814 2379 11878
rect 2443 11814 2460 11878
rect 2524 11814 2541 11878
rect 2605 11814 2622 11878
rect 2686 11814 2703 11878
rect 2767 11814 2784 11878
rect 2848 11814 2865 11878
rect 2929 11814 2946 11878
rect 3010 11814 3027 11878
rect 3091 11814 3108 11878
rect 3172 11814 3189 11878
rect 3253 11814 3270 11878
rect 3334 11814 3351 11878
rect 3415 11814 3432 11878
rect 3496 11814 3513 11878
rect 3577 11814 3594 11878
rect 3658 11814 3675 11878
rect 3739 11814 3756 11878
rect 3820 11814 3837 11878
rect 3901 11814 3918 11878
rect 3982 11814 3999 11878
rect 4063 11814 4080 11878
rect 4144 11814 4161 11878
rect 4225 11814 4242 11878
rect 4306 11814 4323 11878
rect 4387 11814 4404 11878
rect 4468 11814 4485 11878
rect 4549 11814 4566 11878
rect 4630 11814 4647 11878
rect 4711 11814 4728 11878
rect 4792 11814 4809 11878
rect 4873 11814 4874 11878
rect 104 11796 4874 11814
rect 104 11732 105 11796
rect 169 11732 187 11796
rect 251 11732 269 11796
rect 333 11732 351 11796
rect 415 11732 433 11796
rect 497 11732 515 11796
rect 579 11732 597 11796
rect 661 11732 678 11796
rect 742 11732 759 11796
rect 823 11732 840 11796
rect 904 11732 921 11796
rect 985 11732 1002 11796
rect 1066 11732 1083 11796
rect 1147 11732 1164 11796
rect 1228 11732 1245 11796
rect 1309 11732 1326 11796
rect 1390 11732 1407 11796
rect 1471 11732 1488 11796
rect 1552 11732 1569 11796
rect 1633 11732 1650 11796
rect 1714 11732 1731 11796
rect 1795 11732 1812 11796
rect 1876 11732 1893 11796
rect 1957 11732 1974 11796
rect 2038 11732 2055 11796
rect 2119 11732 2136 11796
rect 2200 11732 2217 11796
rect 2281 11732 2298 11796
rect 2362 11732 2379 11796
rect 2443 11732 2460 11796
rect 2524 11732 2541 11796
rect 2605 11732 2622 11796
rect 2686 11732 2703 11796
rect 2767 11732 2784 11796
rect 2848 11732 2865 11796
rect 2929 11732 2946 11796
rect 3010 11732 3027 11796
rect 3091 11732 3108 11796
rect 3172 11732 3189 11796
rect 3253 11732 3270 11796
rect 3334 11732 3351 11796
rect 3415 11732 3432 11796
rect 3496 11732 3513 11796
rect 3577 11732 3594 11796
rect 3658 11732 3675 11796
rect 3739 11732 3756 11796
rect 3820 11732 3837 11796
rect 3901 11732 3918 11796
rect 3982 11732 3999 11796
rect 4063 11732 4080 11796
rect 4144 11732 4161 11796
rect 4225 11732 4242 11796
rect 4306 11732 4323 11796
rect 4387 11732 4404 11796
rect 4468 11732 4485 11796
rect 4549 11732 4566 11796
rect 4630 11732 4647 11796
rect 4711 11732 4728 11796
rect 4792 11732 4809 11796
rect 4873 11732 4874 11796
rect 104 11714 4874 11732
rect 104 11650 105 11714
rect 169 11650 187 11714
rect 251 11650 269 11714
rect 333 11650 351 11714
rect 415 11650 433 11714
rect 497 11650 515 11714
rect 579 11650 597 11714
rect 661 11650 678 11714
rect 742 11650 759 11714
rect 823 11650 840 11714
rect 904 11650 921 11714
rect 985 11650 1002 11714
rect 1066 11650 1083 11714
rect 1147 11650 1164 11714
rect 1228 11650 1245 11714
rect 1309 11650 1326 11714
rect 1390 11650 1407 11714
rect 1471 11650 1488 11714
rect 1552 11650 1569 11714
rect 1633 11650 1650 11714
rect 1714 11650 1731 11714
rect 1795 11650 1812 11714
rect 1876 11650 1893 11714
rect 1957 11650 1974 11714
rect 2038 11650 2055 11714
rect 2119 11650 2136 11714
rect 2200 11650 2217 11714
rect 2281 11650 2298 11714
rect 2362 11650 2379 11714
rect 2443 11650 2460 11714
rect 2524 11650 2541 11714
rect 2605 11650 2622 11714
rect 2686 11650 2703 11714
rect 2767 11650 2784 11714
rect 2848 11650 2865 11714
rect 2929 11650 2946 11714
rect 3010 11650 3027 11714
rect 3091 11650 3108 11714
rect 3172 11650 3189 11714
rect 3253 11650 3270 11714
rect 3334 11650 3351 11714
rect 3415 11650 3432 11714
rect 3496 11650 3513 11714
rect 3577 11650 3594 11714
rect 3658 11650 3675 11714
rect 3739 11650 3756 11714
rect 3820 11650 3837 11714
rect 3901 11650 3918 11714
rect 3982 11650 3999 11714
rect 4063 11650 4080 11714
rect 4144 11650 4161 11714
rect 4225 11650 4242 11714
rect 4306 11650 4323 11714
rect 4387 11650 4404 11714
rect 4468 11650 4485 11714
rect 4549 11650 4566 11714
rect 4630 11650 4647 11714
rect 4711 11650 4728 11714
rect 4792 11650 4809 11714
rect 4873 11650 4874 11714
rect 104 11648 4874 11650
rect 10078 12534 14858 12536
rect 10078 12470 10084 12534
rect 10148 12470 10166 12534
rect 10230 12470 10248 12534
rect 10312 12470 10330 12534
rect 10394 12470 10412 12534
rect 10476 12470 10494 12534
rect 10558 12470 10576 12534
rect 10640 12470 10657 12534
rect 10721 12470 10738 12534
rect 10802 12470 10819 12534
rect 10883 12470 10900 12534
rect 10964 12470 10981 12534
rect 11045 12470 11062 12534
rect 11126 12470 11143 12534
rect 11207 12470 11224 12534
rect 11288 12470 11305 12534
rect 11369 12470 11386 12534
rect 11450 12470 11467 12534
rect 11531 12470 11548 12534
rect 11612 12470 11629 12534
rect 11693 12470 11710 12534
rect 11774 12470 11791 12534
rect 11855 12470 11872 12534
rect 11936 12470 11953 12534
rect 12017 12470 12034 12534
rect 12098 12470 12115 12534
rect 12179 12470 12196 12534
rect 12260 12470 12277 12534
rect 12341 12470 12358 12534
rect 12422 12470 12439 12534
rect 12503 12470 12520 12534
rect 12584 12470 12601 12534
rect 12665 12470 12682 12534
rect 12746 12470 12763 12534
rect 12827 12470 12844 12534
rect 12908 12470 12925 12534
rect 12989 12470 13006 12534
rect 13070 12470 13087 12534
rect 13151 12470 13168 12534
rect 13232 12470 13249 12534
rect 13313 12470 13330 12534
rect 13394 12470 13411 12534
rect 13475 12470 13492 12534
rect 13556 12470 13573 12534
rect 13637 12470 13654 12534
rect 13718 12470 13735 12534
rect 13799 12470 13816 12534
rect 13880 12470 13897 12534
rect 13961 12470 13978 12534
rect 14042 12470 14059 12534
rect 14123 12470 14140 12534
rect 14204 12470 14221 12534
rect 14285 12470 14302 12534
rect 14366 12470 14383 12534
rect 14447 12470 14464 12534
rect 14528 12470 14545 12534
rect 14609 12470 14626 12534
rect 14690 12470 14707 12534
rect 14771 12470 14788 12534
rect 14852 12470 14858 12534
rect 10078 12452 14858 12470
rect 10078 12388 10084 12452
rect 10148 12388 10166 12452
rect 10230 12388 10248 12452
rect 10312 12388 10330 12452
rect 10394 12388 10412 12452
rect 10476 12388 10494 12452
rect 10558 12388 10576 12452
rect 10640 12388 10657 12452
rect 10721 12388 10738 12452
rect 10802 12388 10819 12452
rect 10883 12388 10900 12452
rect 10964 12388 10981 12452
rect 11045 12388 11062 12452
rect 11126 12388 11143 12452
rect 11207 12388 11224 12452
rect 11288 12388 11305 12452
rect 11369 12388 11386 12452
rect 11450 12388 11467 12452
rect 11531 12388 11548 12452
rect 11612 12388 11629 12452
rect 11693 12388 11710 12452
rect 11774 12388 11791 12452
rect 11855 12388 11872 12452
rect 11936 12388 11953 12452
rect 12017 12388 12034 12452
rect 12098 12388 12115 12452
rect 12179 12388 12196 12452
rect 12260 12388 12277 12452
rect 12341 12388 12358 12452
rect 12422 12388 12439 12452
rect 12503 12388 12520 12452
rect 12584 12388 12601 12452
rect 12665 12388 12682 12452
rect 12746 12388 12763 12452
rect 12827 12388 12844 12452
rect 12908 12388 12925 12452
rect 12989 12388 13006 12452
rect 13070 12388 13087 12452
rect 13151 12388 13168 12452
rect 13232 12388 13249 12452
rect 13313 12388 13330 12452
rect 13394 12388 13411 12452
rect 13475 12388 13492 12452
rect 13556 12388 13573 12452
rect 13637 12388 13654 12452
rect 13718 12388 13735 12452
rect 13799 12388 13816 12452
rect 13880 12388 13897 12452
rect 13961 12388 13978 12452
rect 14042 12388 14059 12452
rect 14123 12388 14140 12452
rect 14204 12388 14221 12452
rect 14285 12388 14302 12452
rect 14366 12388 14383 12452
rect 14447 12388 14464 12452
rect 14528 12388 14545 12452
rect 14609 12388 14626 12452
rect 14690 12388 14707 12452
rect 14771 12388 14788 12452
rect 14852 12388 14858 12452
rect 10078 12370 14858 12388
rect 10078 12306 10084 12370
rect 10148 12306 10166 12370
rect 10230 12306 10248 12370
rect 10312 12306 10330 12370
rect 10394 12306 10412 12370
rect 10476 12306 10494 12370
rect 10558 12306 10576 12370
rect 10640 12306 10657 12370
rect 10721 12306 10738 12370
rect 10802 12306 10819 12370
rect 10883 12306 10900 12370
rect 10964 12306 10981 12370
rect 11045 12306 11062 12370
rect 11126 12306 11143 12370
rect 11207 12306 11224 12370
rect 11288 12306 11305 12370
rect 11369 12306 11386 12370
rect 11450 12306 11467 12370
rect 11531 12306 11548 12370
rect 11612 12306 11629 12370
rect 11693 12306 11710 12370
rect 11774 12306 11791 12370
rect 11855 12306 11872 12370
rect 11936 12306 11953 12370
rect 12017 12306 12034 12370
rect 12098 12306 12115 12370
rect 12179 12306 12196 12370
rect 12260 12306 12277 12370
rect 12341 12306 12358 12370
rect 12422 12306 12439 12370
rect 12503 12306 12520 12370
rect 12584 12306 12601 12370
rect 12665 12306 12682 12370
rect 12746 12306 12763 12370
rect 12827 12306 12844 12370
rect 12908 12306 12925 12370
rect 12989 12306 13006 12370
rect 13070 12306 13087 12370
rect 13151 12306 13168 12370
rect 13232 12306 13249 12370
rect 13313 12306 13330 12370
rect 13394 12306 13411 12370
rect 13475 12306 13492 12370
rect 13556 12306 13573 12370
rect 13637 12306 13654 12370
rect 13718 12306 13735 12370
rect 13799 12306 13816 12370
rect 13880 12306 13897 12370
rect 13961 12306 13978 12370
rect 14042 12306 14059 12370
rect 14123 12306 14140 12370
rect 14204 12306 14221 12370
rect 14285 12306 14302 12370
rect 14366 12306 14383 12370
rect 14447 12306 14464 12370
rect 14528 12306 14545 12370
rect 14609 12306 14626 12370
rect 14690 12306 14707 12370
rect 14771 12306 14788 12370
rect 14852 12306 14858 12370
rect 10078 12288 14858 12306
rect 10078 12224 10084 12288
rect 10148 12224 10166 12288
rect 10230 12224 10248 12288
rect 10312 12224 10330 12288
rect 10394 12224 10412 12288
rect 10476 12224 10494 12288
rect 10558 12224 10576 12288
rect 10640 12224 10657 12288
rect 10721 12224 10738 12288
rect 10802 12224 10819 12288
rect 10883 12224 10900 12288
rect 10964 12224 10981 12288
rect 11045 12224 11062 12288
rect 11126 12224 11143 12288
rect 11207 12224 11224 12288
rect 11288 12224 11305 12288
rect 11369 12224 11386 12288
rect 11450 12224 11467 12288
rect 11531 12224 11548 12288
rect 11612 12224 11629 12288
rect 11693 12224 11710 12288
rect 11774 12224 11791 12288
rect 11855 12224 11872 12288
rect 11936 12224 11953 12288
rect 12017 12224 12034 12288
rect 12098 12224 12115 12288
rect 12179 12224 12196 12288
rect 12260 12224 12277 12288
rect 12341 12224 12358 12288
rect 12422 12224 12439 12288
rect 12503 12224 12520 12288
rect 12584 12224 12601 12288
rect 12665 12224 12682 12288
rect 12746 12224 12763 12288
rect 12827 12224 12844 12288
rect 12908 12224 12925 12288
rect 12989 12224 13006 12288
rect 13070 12224 13087 12288
rect 13151 12224 13168 12288
rect 13232 12224 13249 12288
rect 13313 12224 13330 12288
rect 13394 12224 13411 12288
rect 13475 12224 13492 12288
rect 13556 12224 13573 12288
rect 13637 12224 13654 12288
rect 13718 12224 13735 12288
rect 13799 12224 13816 12288
rect 13880 12224 13897 12288
rect 13961 12224 13978 12288
rect 14042 12224 14059 12288
rect 14123 12224 14140 12288
rect 14204 12224 14221 12288
rect 14285 12224 14302 12288
rect 14366 12224 14383 12288
rect 14447 12224 14464 12288
rect 14528 12224 14545 12288
rect 14609 12224 14626 12288
rect 14690 12224 14707 12288
rect 14771 12224 14788 12288
rect 14852 12224 14858 12288
rect 10078 12206 14858 12224
rect 10078 12142 10084 12206
rect 10148 12142 10166 12206
rect 10230 12142 10248 12206
rect 10312 12142 10330 12206
rect 10394 12142 10412 12206
rect 10476 12142 10494 12206
rect 10558 12142 10576 12206
rect 10640 12142 10657 12206
rect 10721 12142 10738 12206
rect 10802 12142 10819 12206
rect 10883 12142 10900 12206
rect 10964 12142 10981 12206
rect 11045 12142 11062 12206
rect 11126 12142 11143 12206
rect 11207 12142 11224 12206
rect 11288 12142 11305 12206
rect 11369 12142 11386 12206
rect 11450 12142 11467 12206
rect 11531 12142 11548 12206
rect 11612 12142 11629 12206
rect 11693 12142 11710 12206
rect 11774 12142 11791 12206
rect 11855 12142 11872 12206
rect 11936 12142 11953 12206
rect 12017 12142 12034 12206
rect 12098 12142 12115 12206
rect 12179 12142 12196 12206
rect 12260 12142 12277 12206
rect 12341 12142 12358 12206
rect 12422 12142 12439 12206
rect 12503 12142 12520 12206
rect 12584 12142 12601 12206
rect 12665 12142 12682 12206
rect 12746 12142 12763 12206
rect 12827 12142 12844 12206
rect 12908 12142 12925 12206
rect 12989 12142 13006 12206
rect 13070 12142 13087 12206
rect 13151 12142 13168 12206
rect 13232 12142 13249 12206
rect 13313 12142 13330 12206
rect 13394 12142 13411 12206
rect 13475 12142 13492 12206
rect 13556 12142 13573 12206
rect 13637 12142 13654 12206
rect 13718 12142 13735 12206
rect 13799 12142 13816 12206
rect 13880 12142 13897 12206
rect 13961 12142 13978 12206
rect 14042 12142 14059 12206
rect 14123 12142 14140 12206
rect 14204 12142 14221 12206
rect 14285 12142 14302 12206
rect 14366 12142 14383 12206
rect 14447 12142 14464 12206
rect 14528 12142 14545 12206
rect 14609 12142 14626 12206
rect 14690 12142 14707 12206
rect 14771 12142 14788 12206
rect 14852 12142 14858 12206
rect 10078 12124 14858 12142
rect 10078 12060 10084 12124
rect 10148 12060 10166 12124
rect 10230 12060 10248 12124
rect 10312 12060 10330 12124
rect 10394 12060 10412 12124
rect 10476 12060 10494 12124
rect 10558 12060 10576 12124
rect 10640 12060 10657 12124
rect 10721 12060 10738 12124
rect 10802 12060 10819 12124
rect 10883 12060 10900 12124
rect 10964 12060 10981 12124
rect 11045 12060 11062 12124
rect 11126 12060 11143 12124
rect 11207 12060 11224 12124
rect 11288 12060 11305 12124
rect 11369 12060 11386 12124
rect 11450 12060 11467 12124
rect 11531 12060 11548 12124
rect 11612 12060 11629 12124
rect 11693 12060 11710 12124
rect 11774 12060 11791 12124
rect 11855 12060 11872 12124
rect 11936 12060 11953 12124
rect 12017 12060 12034 12124
rect 12098 12060 12115 12124
rect 12179 12060 12196 12124
rect 12260 12060 12277 12124
rect 12341 12060 12358 12124
rect 12422 12060 12439 12124
rect 12503 12060 12520 12124
rect 12584 12060 12601 12124
rect 12665 12060 12682 12124
rect 12746 12060 12763 12124
rect 12827 12060 12844 12124
rect 12908 12060 12925 12124
rect 12989 12060 13006 12124
rect 13070 12060 13087 12124
rect 13151 12060 13168 12124
rect 13232 12060 13249 12124
rect 13313 12060 13330 12124
rect 13394 12060 13411 12124
rect 13475 12060 13492 12124
rect 13556 12060 13573 12124
rect 13637 12060 13654 12124
rect 13718 12060 13735 12124
rect 13799 12060 13816 12124
rect 13880 12060 13897 12124
rect 13961 12060 13978 12124
rect 14042 12060 14059 12124
rect 14123 12060 14140 12124
rect 14204 12060 14221 12124
rect 14285 12060 14302 12124
rect 14366 12060 14383 12124
rect 14447 12060 14464 12124
rect 14528 12060 14545 12124
rect 14609 12060 14626 12124
rect 14690 12060 14707 12124
rect 14771 12060 14788 12124
rect 14852 12060 14858 12124
rect 10078 12042 14858 12060
rect 10078 11978 10084 12042
rect 10148 11978 10166 12042
rect 10230 11978 10248 12042
rect 10312 11978 10330 12042
rect 10394 11978 10412 12042
rect 10476 11978 10494 12042
rect 10558 11978 10576 12042
rect 10640 11978 10657 12042
rect 10721 11978 10738 12042
rect 10802 11978 10819 12042
rect 10883 11978 10900 12042
rect 10964 11978 10981 12042
rect 11045 11978 11062 12042
rect 11126 11978 11143 12042
rect 11207 11978 11224 12042
rect 11288 11978 11305 12042
rect 11369 11978 11386 12042
rect 11450 11978 11467 12042
rect 11531 11978 11548 12042
rect 11612 11978 11629 12042
rect 11693 11978 11710 12042
rect 11774 11978 11791 12042
rect 11855 11978 11872 12042
rect 11936 11978 11953 12042
rect 12017 11978 12034 12042
rect 12098 11978 12115 12042
rect 12179 11978 12196 12042
rect 12260 11978 12277 12042
rect 12341 11978 12358 12042
rect 12422 11978 12439 12042
rect 12503 11978 12520 12042
rect 12584 11978 12601 12042
rect 12665 11978 12682 12042
rect 12746 11978 12763 12042
rect 12827 11978 12844 12042
rect 12908 11978 12925 12042
rect 12989 11978 13006 12042
rect 13070 11978 13087 12042
rect 13151 11978 13168 12042
rect 13232 11978 13249 12042
rect 13313 11978 13330 12042
rect 13394 11978 13411 12042
rect 13475 11978 13492 12042
rect 13556 11978 13573 12042
rect 13637 11978 13654 12042
rect 13718 11978 13735 12042
rect 13799 11978 13816 12042
rect 13880 11978 13897 12042
rect 13961 11978 13978 12042
rect 14042 11978 14059 12042
rect 14123 11978 14140 12042
rect 14204 11978 14221 12042
rect 14285 11978 14302 12042
rect 14366 11978 14383 12042
rect 14447 11978 14464 12042
rect 14528 11978 14545 12042
rect 14609 11978 14626 12042
rect 14690 11978 14707 12042
rect 14771 11978 14788 12042
rect 14852 11978 14858 12042
rect 10078 11960 14858 11978
rect 10078 11896 10084 11960
rect 10148 11896 10166 11960
rect 10230 11896 10248 11960
rect 10312 11896 10330 11960
rect 10394 11896 10412 11960
rect 10476 11896 10494 11960
rect 10558 11896 10576 11960
rect 10640 11896 10657 11960
rect 10721 11896 10738 11960
rect 10802 11896 10819 11960
rect 10883 11896 10900 11960
rect 10964 11896 10981 11960
rect 11045 11896 11062 11960
rect 11126 11896 11143 11960
rect 11207 11896 11224 11960
rect 11288 11896 11305 11960
rect 11369 11896 11386 11960
rect 11450 11896 11467 11960
rect 11531 11896 11548 11960
rect 11612 11896 11629 11960
rect 11693 11896 11710 11960
rect 11774 11896 11791 11960
rect 11855 11896 11872 11960
rect 11936 11896 11953 11960
rect 12017 11896 12034 11960
rect 12098 11896 12115 11960
rect 12179 11896 12196 11960
rect 12260 11896 12277 11960
rect 12341 11896 12358 11960
rect 12422 11896 12439 11960
rect 12503 11896 12520 11960
rect 12584 11896 12601 11960
rect 12665 11896 12682 11960
rect 12746 11896 12763 11960
rect 12827 11896 12844 11960
rect 12908 11896 12925 11960
rect 12989 11896 13006 11960
rect 13070 11896 13087 11960
rect 13151 11896 13168 11960
rect 13232 11896 13249 11960
rect 13313 11896 13330 11960
rect 13394 11896 13411 11960
rect 13475 11896 13492 11960
rect 13556 11896 13573 11960
rect 13637 11896 13654 11960
rect 13718 11896 13735 11960
rect 13799 11896 13816 11960
rect 13880 11896 13897 11960
rect 13961 11896 13978 11960
rect 14042 11896 14059 11960
rect 14123 11896 14140 11960
rect 14204 11896 14221 11960
rect 14285 11896 14302 11960
rect 14366 11896 14383 11960
rect 14447 11896 14464 11960
rect 14528 11896 14545 11960
rect 14609 11896 14626 11960
rect 14690 11896 14707 11960
rect 14771 11896 14788 11960
rect 14852 11896 14858 11960
rect 10078 11878 14858 11896
rect 10078 11814 10084 11878
rect 10148 11814 10166 11878
rect 10230 11814 10248 11878
rect 10312 11814 10330 11878
rect 10394 11814 10412 11878
rect 10476 11814 10494 11878
rect 10558 11814 10576 11878
rect 10640 11814 10657 11878
rect 10721 11814 10738 11878
rect 10802 11814 10819 11878
rect 10883 11814 10900 11878
rect 10964 11814 10981 11878
rect 11045 11814 11062 11878
rect 11126 11814 11143 11878
rect 11207 11814 11224 11878
rect 11288 11814 11305 11878
rect 11369 11814 11386 11878
rect 11450 11814 11467 11878
rect 11531 11814 11548 11878
rect 11612 11814 11629 11878
rect 11693 11814 11710 11878
rect 11774 11814 11791 11878
rect 11855 11814 11872 11878
rect 11936 11814 11953 11878
rect 12017 11814 12034 11878
rect 12098 11814 12115 11878
rect 12179 11814 12196 11878
rect 12260 11814 12277 11878
rect 12341 11814 12358 11878
rect 12422 11814 12439 11878
rect 12503 11814 12520 11878
rect 12584 11814 12601 11878
rect 12665 11814 12682 11878
rect 12746 11814 12763 11878
rect 12827 11814 12844 11878
rect 12908 11814 12925 11878
rect 12989 11814 13006 11878
rect 13070 11814 13087 11878
rect 13151 11814 13168 11878
rect 13232 11814 13249 11878
rect 13313 11814 13330 11878
rect 13394 11814 13411 11878
rect 13475 11814 13492 11878
rect 13556 11814 13573 11878
rect 13637 11814 13654 11878
rect 13718 11814 13735 11878
rect 13799 11814 13816 11878
rect 13880 11814 13897 11878
rect 13961 11814 13978 11878
rect 14042 11814 14059 11878
rect 14123 11814 14140 11878
rect 14204 11814 14221 11878
rect 14285 11814 14302 11878
rect 14366 11814 14383 11878
rect 14447 11814 14464 11878
rect 14528 11814 14545 11878
rect 14609 11814 14626 11878
rect 14690 11814 14707 11878
rect 14771 11814 14788 11878
rect 14852 11814 14858 11878
rect 10078 11796 14858 11814
rect 10078 11732 10084 11796
rect 10148 11732 10166 11796
rect 10230 11732 10248 11796
rect 10312 11732 10330 11796
rect 10394 11732 10412 11796
rect 10476 11732 10494 11796
rect 10558 11732 10576 11796
rect 10640 11732 10657 11796
rect 10721 11732 10738 11796
rect 10802 11732 10819 11796
rect 10883 11732 10900 11796
rect 10964 11732 10981 11796
rect 11045 11732 11062 11796
rect 11126 11732 11143 11796
rect 11207 11732 11224 11796
rect 11288 11732 11305 11796
rect 11369 11732 11386 11796
rect 11450 11732 11467 11796
rect 11531 11732 11548 11796
rect 11612 11732 11629 11796
rect 11693 11732 11710 11796
rect 11774 11732 11791 11796
rect 11855 11732 11872 11796
rect 11936 11732 11953 11796
rect 12017 11732 12034 11796
rect 12098 11732 12115 11796
rect 12179 11732 12196 11796
rect 12260 11732 12277 11796
rect 12341 11732 12358 11796
rect 12422 11732 12439 11796
rect 12503 11732 12520 11796
rect 12584 11732 12601 11796
rect 12665 11732 12682 11796
rect 12746 11732 12763 11796
rect 12827 11732 12844 11796
rect 12908 11732 12925 11796
rect 12989 11732 13006 11796
rect 13070 11732 13087 11796
rect 13151 11732 13168 11796
rect 13232 11732 13249 11796
rect 13313 11732 13330 11796
rect 13394 11732 13411 11796
rect 13475 11732 13492 11796
rect 13556 11732 13573 11796
rect 13637 11732 13654 11796
rect 13718 11732 13735 11796
rect 13799 11732 13816 11796
rect 13880 11732 13897 11796
rect 13961 11732 13978 11796
rect 14042 11732 14059 11796
rect 14123 11732 14140 11796
rect 14204 11732 14221 11796
rect 14285 11732 14302 11796
rect 14366 11732 14383 11796
rect 14447 11732 14464 11796
rect 14528 11732 14545 11796
rect 14609 11732 14626 11796
rect 14690 11732 14707 11796
rect 14771 11732 14788 11796
rect 14852 11732 14858 11796
rect 10078 11714 14858 11732
rect 10078 11650 10084 11714
rect 10148 11650 10166 11714
rect 10230 11650 10248 11714
rect 10312 11650 10330 11714
rect 10394 11650 10412 11714
rect 10476 11650 10494 11714
rect 10558 11650 10576 11714
rect 10640 11650 10657 11714
rect 10721 11650 10738 11714
rect 10802 11650 10819 11714
rect 10883 11650 10900 11714
rect 10964 11650 10981 11714
rect 11045 11650 11062 11714
rect 11126 11650 11143 11714
rect 11207 11650 11224 11714
rect 11288 11650 11305 11714
rect 11369 11650 11386 11714
rect 11450 11650 11467 11714
rect 11531 11650 11548 11714
rect 11612 11650 11629 11714
rect 11693 11650 11710 11714
rect 11774 11650 11791 11714
rect 11855 11650 11872 11714
rect 11936 11650 11953 11714
rect 12017 11650 12034 11714
rect 12098 11650 12115 11714
rect 12179 11650 12196 11714
rect 12260 11650 12277 11714
rect 12341 11650 12358 11714
rect 12422 11650 12439 11714
rect 12503 11650 12520 11714
rect 12584 11650 12601 11714
rect 12665 11650 12682 11714
rect 12746 11650 12763 11714
rect 12827 11650 12844 11714
rect 12908 11650 12925 11714
rect 12989 11650 13006 11714
rect 13070 11650 13087 11714
rect 13151 11650 13168 11714
rect 13232 11650 13249 11714
rect 13313 11650 13330 11714
rect 13394 11650 13411 11714
rect 13475 11650 13492 11714
rect 13556 11650 13573 11714
rect 13637 11650 13654 11714
rect 13718 11650 13735 11714
rect 13799 11650 13816 11714
rect 13880 11650 13897 11714
rect 13961 11650 13978 11714
rect 14042 11650 14059 11714
rect 14123 11650 14140 11714
rect 14204 11650 14221 11714
rect 14285 11650 14302 11714
rect 14366 11650 14383 11714
rect 14447 11650 14464 11714
rect 14528 11650 14545 11714
rect 14609 11650 14626 11714
rect 14690 11650 14707 11714
rect 14771 11650 14788 11714
rect 14852 11650 14858 11714
rect 10078 11648 14858 11650
rect 99 6094 4879 6096
rect 99 6030 105 6094
rect 169 6030 187 6094
rect 251 6030 269 6094
rect 333 6030 351 6094
rect 415 6030 433 6094
rect 497 6030 515 6094
rect 579 6030 597 6094
rect 661 6030 678 6094
rect 742 6030 759 6094
rect 823 6030 840 6094
rect 904 6030 921 6094
rect 985 6030 1002 6094
rect 1066 6030 1083 6094
rect 1147 6030 1164 6094
rect 1228 6030 1245 6094
rect 1309 6030 1326 6094
rect 1390 6030 1407 6094
rect 1471 6030 1488 6094
rect 1552 6030 1569 6094
rect 1633 6030 1650 6094
rect 1714 6030 1731 6094
rect 1795 6030 1812 6094
rect 1876 6030 1893 6094
rect 1957 6030 1974 6094
rect 2038 6030 2055 6094
rect 2119 6030 2136 6094
rect 2200 6030 2217 6094
rect 2281 6030 2298 6094
rect 2362 6030 2379 6094
rect 2443 6030 2460 6094
rect 2524 6030 2541 6094
rect 2605 6030 2622 6094
rect 2686 6030 2703 6094
rect 2767 6030 2784 6094
rect 2848 6030 2865 6094
rect 2929 6030 2946 6094
rect 3010 6030 3027 6094
rect 3091 6030 3108 6094
rect 3172 6030 3189 6094
rect 3253 6030 3270 6094
rect 3334 6030 3351 6094
rect 3415 6030 3432 6094
rect 3496 6030 3513 6094
rect 3577 6030 3594 6094
rect 3658 6030 3675 6094
rect 3739 6030 3756 6094
rect 3820 6030 3837 6094
rect 3901 6030 3918 6094
rect 3982 6030 3999 6094
rect 4063 6030 4080 6094
rect 4144 6030 4161 6094
rect 4225 6030 4242 6094
rect 4306 6030 4323 6094
rect 4387 6030 4404 6094
rect 4468 6030 4485 6094
rect 4549 6030 4566 6094
rect 4630 6030 4647 6094
rect 4711 6030 4728 6094
rect 4792 6030 4809 6094
rect 4873 6030 4879 6094
rect 99 6008 4879 6030
rect 99 5944 105 6008
rect 169 5944 187 6008
rect 251 5944 269 6008
rect 333 5944 351 6008
rect 415 5944 433 6008
rect 497 5944 515 6008
rect 579 5944 597 6008
rect 661 5944 678 6008
rect 742 5944 759 6008
rect 823 5944 840 6008
rect 904 5944 921 6008
rect 985 5944 1002 6008
rect 1066 5944 1083 6008
rect 1147 5944 1164 6008
rect 1228 5944 1245 6008
rect 1309 5944 1326 6008
rect 1390 5944 1407 6008
rect 1471 5944 1488 6008
rect 1552 5944 1569 6008
rect 1633 5944 1650 6008
rect 1714 5944 1731 6008
rect 1795 5944 1812 6008
rect 1876 5944 1893 6008
rect 1957 5944 1974 6008
rect 2038 5944 2055 6008
rect 2119 5944 2136 6008
rect 2200 5944 2217 6008
rect 2281 5944 2298 6008
rect 2362 5944 2379 6008
rect 2443 5944 2460 6008
rect 2524 5944 2541 6008
rect 2605 5944 2622 6008
rect 2686 5944 2703 6008
rect 2767 5944 2784 6008
rect 2848 5944 2865 6008
rect 2929 5944 2946 6008
rect 3010 5944 3027 6008
rect 3091 5944 3108 6008
rect 3172 5944 3189 6008
rect 3253 5944 3270 6008
rect 3334 5944 3351 6008
rect 3415 5944 3432 6008
rect 3496 5944 3513 6008
rect 3577 5944 3594 6008
rect 3658 5944 3675 6008
rect 3739 5944 3756 6008
rect 3820 5944 3837 6008
rect 3901 5944 3918 6008
rect 3982 5944 3999 6008
rect 4063 5944 4080 6008
rect 4144 5944 4161 6008
rect 4225 5944 4242 6008
rect 4306 5944 4323 6008
rect 4387 5944 4404 6008
rect 4468 5944 4485 6008
rect 4549 5944 4566 6008
rect 4630 5944 4647 6008
rect 4711 5944 4728 6008
rect 4792 5944 4809 6008
rect 4873 5944 4879 6008
rect 99 5922 4879 5944
rect 99 5858 105 5922
rect 169 5858 187 5922
rect 251 5858 269 5922
rect 333 5858 351 5922
rect 415 5858 433 5922
rect 497 5858 515 5922
rect 579 5858 597 5922
rect 661 5858 678 5922
rect 742 5858 759 5922
rect 823 5858 840 5922
rect 904 5858 921 5922
rect 985 5858 1002 5922
rect 1066 5858 1083 5922
rect 1147 5858 1164 5922
rect 1228 5858 1245 5922
rect 1309 5858 1326 5922
rect 1390 5858 1407 5922
rect 1471 5858 1488 5922
rect 1552 5858 1569 5922
rect 1633 5858 1650 5922
rect 1714 5858 1731 5922
rect 1795 5858 1812 5922
rect 1876 5858 1893 5922
rect 1957 5858 1974 5922
rect 2038 5858 2055 5922
rect 2119 5858 2136 5922
rect 2200 5858 2217 5922
rect 2281 5858 2298 5922
rect 2362 5858 2379 5922
rect 2443 5858 2460 5922
rect 2524 5858 2541 5922
rect 2605 5858 2622 5922
rect 2686 5858 2703 5922
rect 2767 5858 2784 5922
rect 2848 5858 2865 5922
rect 2929 5858 2946 5922
rect 3010 5858 3027 5922
rect 3091 5858 3108 5922
rect 3172 5858 3189 5922
rect 3253 5858 3270 5922
rect 3334 5858 3351 5922
rect 3415 5858 3432 5922
rect 3496 5858 3513 5922
rect 3577 5858 3594 5922
rect 3658 5858 3675 5922
rect 3739 5858 3756 5922
rect 3820 5858 3837 5922
rect 3901 5858 3918 5922
rect 3982 5858 3999 5922
rect 4063 5858 4080 5922
rect 4144 5858 4161 5922
rect 4225 5858 4242 5922
rect 4306 5858 4323 5922
rect 4387 5858 4404 5922
rect 4468 5858 4485 5922
rect 4549 5858 4566 5922
rect 4630 5858 4647 5922
rect 4711 5858 4728 5922
rect 4792 5858 4809 5922
rect 4873 5858 4879 5922
rect 99 5836 4879 5858
rect 99 5772 105 5836
rect 169 5772 187 5836
rect 251 5772 269 5836
rect 333 5772 351 5836
rect 415 5772 433 5836
rect 497 5772 515 5836
rect 579 5772 597 5836
rect 661 5772 678 5836
rect 742 5772 759 5836
rect 823 5772 840 5836
rect 904 5772 921 5836
rect 985 5772 1002 5836
rect 1066 5772 1083 5836
rect 1147 5772 1164 5836
rect 1228 5772 1245 5836
rect 1309 5772 1326 5836
rect 1390 5772 1407 5836
rect 1471 5772 1488 5836
rect 1552 5772 1569 5836
rect 1633 5772 1650 5836
rect 1714 5772 1731 5836
rect 1795 5772 1812 5836
rect 1876 5772 1893 5836
rect 1957 5772 1974 5836
rect 2038 5772 2055 5836
rect 2119 5772 2136 5836
rect 2200 5772 2217 5836
rect 2281 5772 2298 5836
rect 2362 5772 2379 5836
rect 2443 5772 2460 5836
rect 2524 5772 2541 5836
rect 2605 5772 2622 5836
rect 2686 5772 2703 5836
rect 2767 5772 2784 5836
rect 2848 5772 2865 5836
rect 2929 5772 2946 5836
rect 3010 5772 3027 5836
rect 3091 5772 3108 5836
rect 3172 5772 3189 5836
rect 3253 5772 3270 5836
rect 3334 5772 3351 5836
rect 3415 5772 3432 5836
rect 3496 5772 3513 5836
rect 3577 5772 3594 5836
rect 3658 5772 3675 5836
rect 3739 5772 3756 5836
rect 3820 5772 3837 5836
rect 3901 5772 3918 5836
rect 3982 5772 3999 5836
rect 4063 5772 4080 5836
rect 4144 5772 4161 5836
rect 4225 5772 4242 5836
rect 4306 5772 4323 5836
rect 4387 5772 4404 5836
rect 4468 5772 4485 5836
rect 4549 5772 4566 5836
rect 4630 5772 4647 5836
rect 4711 5772 4728 5836
rect 4792 5772 4809 5836
rect 4873 5772 4879 5836
rect 99 5750 4879 5772
rect 99 5686 105 5750
rect 169 5686 187 5750
rect 251 5686 269 5750
rect 333 5686 351 5750
rect 415 5686 433 5750
rect 497 5686 515 5750
rect 579 5686 597 5750
rect 661 5686 678 5750
rect 742 5686 759 5750
rect 823 5686 840 5750
rect 904 5686 921 5750
rect 985 5686 1002 5750
rect 1066 5686 1083 5750
rect 1147 5686 1164 5750
rect 1228 5686 1245 5750
rect 1309 5686 1326 5750
rect 1390 5686 1407 5750
rect 1471 5686 1488 5750
rect 1552 5686 1569 5750
rect 1633 5686 1650 5750
rect 1714 5686 1731 5750
rect 1795 5686 1812 5750
rect 1876 5686 1893 5750
rect 1957 5686 1974 5750
rect 2038 5686 2055 5750
rect 2119 5686 2136 5750
rect 2200 5686 2217 5750
rect 2281 5686 2298 5750
rect 2362 5686 2379 5750
rect 2443 5686 2460 5750
rect 2524 5686 2541 5750
rect 2605 5686 2622 5750
rect 2686 5686 2703 5750
rect 2767 5686 2784 5750
rect 2848 5686 2865 5750
rect 2929 5686 2946 5750
rect 3010 5686 3027 5750
rect 3091 5686 3108 5750
rect 3172 5686 3189 5750
rect 3253 5686 3270 5750
rect 3334 5686 3351 5750
rect 3415 5686 3432 5750
rect 3496 5686 3513 5750
rect 3577 5686 3594 5750
rect 3658 5686 3675 5750
rect 3739 5686 3756 5750
rect 3820 5686 3837 5750
rect 3901 5686 3918 5750
rect 3982 5686 3999 5750
rect 4063 5686 4080 5750
rect 4144 5686 4161 5750
rect 4225 5686 4242 5750
rect 4306 5686 4323 5750
rect 4387 5686 4404 5750
rect 4468 5686 4485 5750
rect 4549 5686 4566 5750
rect 4630 5686 4647 5750
rect 4711 5686 4728 5750
rect 4792 5686 4809 5750
rect 4873 5686 4879 5750
rect 99 5664 4879 5686
rect 99 5600 105 5664
rect 169 5600 187 5664
rect 251 5600 269 5664
rect 333 5600 351 5664
rect 415 5600 433 5664
rect 497 5600 515 5664
rect 579 5600 597 5664
rect 661 5600 678 5664
rect 742 5600 759 5664
rect 823 5600 840 5664
rect 904 5600 921 5664
rect 985 5600 1002 5664
rect 1066 5600 1083 5664
rect 1147 5600 1164 5664
rect 1228 5600 1245 5664
rect 1309 5600 1326 5664
rect 1390 5600 1407 5664
rect 1471 5600 1488 5664
rect 1552 5600 1569 5664
rect 1633 5600 1650 5664
rect 1714 5600 1731 5664
rect 1795 5600 1812 5664
rect 1876 5600 1893 5664
rect 1957 5600 1974 5664
rect 2038 5600 2055 5664
rect 2119 5600 2136 5664
rect 2200 5600 2217 5664
rect 2281 5600 2298 5664
rect 2362 5600 2379 5664
rect 2443 5600 2460 5664
rect 2524 5600 2541 5664
rect 2605 5600 2622 5664
rect 2686 5600 2703 5664
rect 2767 5600 2784 5664
rect 2848 5600 2865 5664
rect 2929 5600 2946 5664
rect 3010 5600 3027 5664
rect 3091 5600 3108 5664
rect 3172 5600 3189 5664
rect 3253 5600 3270 5664
rect 3334 5600 3351 5664
rect 3415 5600 3432 5664
rect 3496 5600 3513 5664
rect 3577 5600 3594 5664
rect 3658 5600 3675 5664
rect 3739 5600 3756 5664
rect 3820 5600 3837 5664
rect 3901 5600 3918 5664
rect 3982 5600 3999 5664
rect 4063 5600 4080 5664
rect 4144 5600 4161 5664
rect 4225 5600 4242 5664
rect 4306 5600 4323 5664
rect 4387 5600 4404 5664
rect 4468 5600 4485 5664
rect 4549 5600 4566 5664
rect 4630 5600 4647 5664
rect 4711 5600 4728 5664
rect 4792 5600 4809 5664
rect 4873 5600 4879 5664
rect 99 5578 4879 5600
rect 99 5514 105 5578
rect 169 5514 187 5578
rect 251 5514 269 5578
rect 333 5514 351 5578
rect 415 5514 433 5578
rect 497 5514 515 5578
rect 579 5514 597 5578
rect 661 5514 678 5578
rect 742 5514 759 5578
rect 823 5514 840 5578
rect 904 5514 921 5578
rect 985 5514 1002 5578
rect 1066 5514 1083 5578
rect 1147 5514 1164 5578
rect 1228 5514 1245 5578
rect 1309 5514 1326 5578
rect 1390 5514 1407 5578
rect 1471 5514 1488 5578
rect 1552 5514 1569 5578
rect 1633 5514 1650 5578
rect 1714 5514 1731 5578
rect 1795 5514 1812 5578
rect 1876 5514 1893 5578
rect 1957 5514 1974 5578
rect 2038 5514 2055 5578
rect 2119 5514 2136 5578
rect 2200 5514 2217 5578
rect 2281 5514 2298 5578
rect 2362 5514 2379 5578
rect 2443 5514 2460 5578
rect 2524 5514 2541 5578
rect 2605 5514 2622 5578
rect 2686 5514 2703 5578
rect 2767 5514 2784 5578
rect 2848 5514 2865 5578
rect 2929 5514 2946 5578
rect 3010 5514 3027 5578
rect 3091 5514 3108 5578
rect 3172 5514 3189 5578
rect 3253 5514 3270 5578
rect 3334 5514 3351 5578
rect 3415 5514 3432 5578
rect 3496 5514 3513 5578
rect 3577 5514 3594 5578
rect 3658 5514 3675 5578
rect 3739 5514 3756 5578
rect 3820 5514 3837 5578
rect 3901 5514 3918 5578
rect 3982 5514 3999 5578
rect 4063 5514 4080 5578
rect 4144 5514 4161 5578
rect 4225 5514 4242 5578
rect 4306 5514 4323 5578
rect 4387 5514 4404 5578
rect 4468 5514 4485 5578
rect 4549 5514 4566 5578
rect 4630 5514 4647 5578
rect 4711 5514 4728 5578
rect 4792 5514 4809 5578
rect 4873 5514 4879 5578
rect 99 5492 4879 5514
rect 99 5428 105 5492
rect 169 5428 187 5492
rect 251 5428 269 5492
rect 333 5428 351 5492
rect 415 5428 433 5492
rect 497 5428 515 5492
rect 579 5428 597 5492
rect 661 5428 678 5492
rect 742 5428 759 5492
rect 823 5428 840 5492
rect 904 5428 921 5492
rect 985 5428 1002 5492
rect 1066 5428 1083 5492
rect 1147 5428 1164 5492
rect 1228 5428 1245 5492
rect 1309 5428 1326 5492
rect 1390 5428 1407 5492
rect 1471 5428 1488 5492
rect 1552 5428 1569 5492
rect 1633 5428 1650 5492
rect 1714 5428 1731 5492
rect 1795 5428 1812 5492
rect 1876 5428 1893 5492
rect 1957 5428 1974 5492
rect 2038 5428 2055 5492
rect 2119 5428 2136 5492
rect 2200 5428 2217 5492
rect 2281 5428 2298 5492
rect 2362 5428 2379 5492
rect 2443 5428 2460 5492
rect 2524 5428 2541 5492
rect 2605 5428 2622 5492
rect 2686 5428 2703 5492
rect 2767 5428 2784 5492
rect 2848 5428 2865 5492
rect 2929 5428 2946 5492
rect 3010 5428 3027 5492
rect 3091 5428 3108 5492
rect 3172 5428 3189 5492
rect 3253 5428 3270 5492
rect 3334 5428 3351 5492
rect 3415 5428 3432 5492
rect 3496 5428 3513 5492
rect 3577 5428 3594 5492
rect 3658 5428 3675 5492
rect 3739 5428 3756 5492
rect 3820 5428 3837 5492
rect 3901 5428 3918 5492
rect 3982 5428 3999 5492
rect 4063 5428 4080 5492
rect 4144 5428 4161 5492
rect 4225 5428 4242 5492
rect 4306 5428 4323 5492
rect 4387 5428 4404 5492
rect 4468 5428 4485 5492
rect 4549 5428 4566 5492
rect 4630 5428 4647 5492
rect 4711 5428 4728 5492
rect 4792 5428 4809 5492
rect 4873 5428 4879 5492
rect 99 5406 4879 5428
rect 99 5342 105 5406
rect 169 5342 187 5406
rect 251 5342 269 5406
rect 333 5342 351 5406
rect 415 5342 433 5406
rect 497 5342 515 5406
rect 579 5342 597 5406
rect 661 5342 678 5406
rect 742 5342 759 5406
rect 823 5342 840 5406
rect 904 5342 921 5406
rect 985 5342 1002 5406
rect 1066 5342 1083 5406
rect 1147 5342 1164 5406
rect 1228 5342 1245 5406
rect 1309 5342 1326 5406
rect 1390 5342 1407 5406
rect 1471 5342 1488 5406
rect 1552 5342 1569 5406
rect 1633 5342 1650 5406
rect 1714 5342 1731 5406
rect 1795 5342 1812 5406
rect 1876 5342 1893 5406
rect 1957 5342 1974 5406
rect 2038 5342 2055 5406
rect 2119 5342 2136 5406
rect 2200 5342 2217 5406
rect 2281 5342 2298 5406
rect 2362 5342 2379 5406
rect 2443 5342 2460 5406
rect 2524 5342 2541 5406
rect 2605 5342 2622 5406
rect 2686 5342 2703 5406
rect 2767 5342 2784 5406
rect 2848 5342 2865 5406
rect 2929 5342 2946 5406
rect 3010 5342 3027 5406
rect 3091 5342 3108 5406
rect 3172 5342 3189 5406
rect 3253 5342 3270 5406
rect 3334 5342 3351 5406
rect 3415 5342 3432 5406
rect 3496 5342 3513 5406
rect 3577 5342 3594 5406
rect 3658 5342 3675 5406
rect 3739 5342 3756 5406
rect 3820 5342 3837 5406
rect 3901 5342 3918 5406
rect 3982 5342 3999 5406
rect 4063 5342 4080 5406
rect 4144 5342 4161 5406
rect 4225 5342 4242 5406
rect 4306 5342 4323 5406
rect 4387 5342 4404 5406
rect 4468 5342 4485 5406
rect 4549 5342 4566 5406
rect 4630 5342 4647 5406
rect 4711 5342 4728 5406
rect 4792 5342 4809 5406
rect 4873 5342 4879 5406
rect 99 5320 4879 5342
rect 99 5256 105 5320
rect 169 5256 187 5320
rect 251 5256 269 5320
rect 333 5256 351 5320
rect 415 5256 433 5320
rect 497 5256 515 5320
rect 579 5256 597 5320
rect 661 5256 678 5320
rect 742 5256 759 5320
rect 823 5256 840 5320
rect 904 5256 921 5320
rect 985 5256 1002 5320
rect 1066 5256 1083 5320
rect 1147 5256 1164 5320
rect 1228 5256 1245 5320
rect 1309 5256 1326 5320
rect 1390 5256 1407 5320
rect 1471 5256 1488 5320
rect 1552 5256 1569 5320
rect 1633 5256 1650 5320
rect 1714 5256 1731 5320
rect 1795 5256 1812 5320
rect 1876 5256 1893 5320
rect 1957 5256 1974 5320
rect 2038 5256 2055 5320
rect 2119 5256 2136 5320
rect 2200 5256 2217 5320
rect 2281 5256 2298 5320
rect 2362 5256 2379 5320
rect 2443 5256 2460 5320
rect 2524 5256 2541 5320
rect 2605 5256 2622 5320
rect 2686 5256 2703 5320
rect 2767 5256 2784 5320
rect 2848 5256 2865 5320
rect 2929 5256 2946 5320
rect 3010 5256 3027 5320
rect 3091 5256 3108 5320
rect 3172 5256 3189 5320
rect 3253 5256 3270 5320
rect 3334 5256 3351 5320
rect 3415 5256 3432 5320
rect 3496 5256 3513 5320
rect 3577 5256 3594 5320
rect 3658 5256 3675 5320
rect 3739 5256 3756 5320
rect 3820 5256 3837 5320
rect 3901 5256 3918 5320
rect 3982 5256 3999 5320
rect 4063 5256 4080 5320
rect 4144 5256 4161 5320
rect 4225 5256 4242 5320
rect 4306 5256 4323 5320
rect 4387 5256 4404 5320
rect 4468 5256 4485 5320
rect 4549 5256 4566 5320
rect 4630 5256 4647 5320
rect 4711 5256 4728 5320
rect 4792 5256 4809 5320
rect 4873 5256 4879 5320
rect 99 5234 4879 5256
rect 99 5170 105 5234
rect 169 5170 187 5234
rect 251 5170 269 5234
rect 333 5170 351 5234
rect 415 5170 433 5234
rect 497 5170 515 5234
rect 579 5170 597 5234
rect 661 5170 678 5234
rect 742 5170 759 5234
rect 823 5170 840 5234
rect 904 5170 921 5234
rect 985 5170 1002 5234
rect 1066 5170 1083 5234
rect 1147 5170 1164 5234
rect 1228 5170 1245 5234
rect 1309 5170 1326 5234
rect 1390 5170 1407 5234
rect 1471 5170 1488 5234
rect 1552 5170 1569 5234
rect 1633 5170 1650 5234
rect 1714 5170 1731 5234
rect 1795 5170 1812 5234
rect 1876 5170 1893 5234
rect 1957 5170 1974 5234
rect 2038 5170 2055 5234
rect 2119 5170 2136 5234
rect 2200 5170 2217 5234
rect 2281 5170 2298 5234
rect 2362 5170 2379 5234
rect 2443 5170 2460 5234
rect 2524 5170 2541 5234
rect 2605 5170 2622 5234
rect 2686 5170 2703 5234
rect 2767 5170 2784 5234
rect 2848 5170 2865 5234
rect 2929 5170 2946 5234
rect 3010 5170 3027 5234
rect 3091 5170 3108 5234
rect 3172 5170 3189 5234
rect 3253 5170 3270 5234
rect 3334 5170 3351 5234
rect 3415 5170 3432 5234
rect 3496 5170 3513 5234
rect 3577 5170 3594 5234
rect 3658 5170 3675 5234
rect 3739 5170 3756 5234
rect 3820 5170 3837 5234
rect 3901 5170 3918 5234
rect 3982 5170 3999 5234
rect 4063 5170 4080 5234
rect 4144 5170 4161 5234
rect 4225 5170 4242 5234
rect 4306 5170 4323 5234
rect 4387 5170 4404 5234
rect 4468 5170 4485 5234
rect 4549 5170 4566 5234
rect 4630 5170 4647 5234
rect 4711 5170 4728 5234
rect 4792 5170 4809 5234
rect 4873 5170 4879 5234
rect 99 5168 4879 5170
rect 10078 6094 14858 6096
rect 10078 6030 10084 6094
rect 10148 6030 10166 6094
rect 10230 6030 10248 6094
rect 10312 6030 10330 6094
rect 10394 6030 10412 6094
rect 10476 6030 10494 6094
rect 10558 6030 10576 6094
rect 10640 6030 10657 6094
rect 10721 6030 10738 6094
rect 10802 6030 10819 6094
rect 10883 6030 10900 6094
rect 10964 6030 10981 6094
rect 11045 6030 11062 6094
rect 11126 6030 11143 6094
rect 11207 6030 11224 6094
rect 11288 6030 11305 6094
rect 11369 6030 11386 6094
rect 11450 6030 11467 6094
rect 11531 6030 11548 6094
rect 11612 6030 11629 6094
rect 11693 6030 11710 6094
rect 11774 6030 11791 6094
rect 11855 6030 11872 6094
rect 11936 6030 11953 6094
rect 12017 6030 12034 6094
rect 12098 6030 12115 6094
rect 12179 6030 12196 6094
rect 12260 6030 12277 6094
rect 12341 6030 12358 6094
rect 12422 6030 12439 6094
rect 12503 6030 12520 6094
rect 12584 6030 12601 6094
rect 12665 6030 12682 6094
rect 12746 6030 12763 6094
rect 12827 6030 12844 6094
rect 12908 6030 12925 6094
rect 12989 6030 13006 6094
rect 13070 6030 13087 6094
rect 13151 6030 13168 6094
rect 13232 6030 13249 6094
rect 13313 6030 13330 6094
rect 13394 6030 13411 6094
rect 13475 6030 13492 6094
rect 13556 6030 13573 6094
rect 13637 6030 13654 6094
rect 13718 6030 13735 6094
rect 13799 6030 13816 6094
rect 13880 6030 13897 6094
rect 13961 6030 13978 6094
rect 14042 6030 14059 6094
rect 14123 6030 14140 6094
rect 14204 6030 14221 6094
rect 14285 6030 14302 6094
rect 14366 6030 14383 6094
rect 14447 6030 14464 6094
rect 14528 6030 14545 6094
rect 14609 6030 14626 6094
rect 14690 6030 14707 6094
rect 14771 6030 14788 6094
rect 14852 6030 14858 6094
rect 10078 6008 14858 6030
rect 10078 5944 10084 6008
rect 10148 5944 10166 6008
rect 10230 5944 10248 6008
rect 10312 5944 10330 6008
rect 10394 5944 10412 6008
rect 10476 5944 10494 6008
rect 10558 5944 10576 6008
rect 10640 5944 10657 6008
rect 10721 5944 10738 6008
rect 10802 5944 10819 6008
rect 10883 5944 10900 6008
rect 10964 5944 10981 6008
rect 11045 5944 11062 6008
rect 11126 5944 11143 6008
rect 11207 5944 11224 6008
rect 11288 5944 11305 6008
rect 11369 5944 11386 6008
rect 11450 5944 11467 6008
rect 11531 5944 11548 6008
rect 11612 5944 11629 6008
rect 11693 5944 11710 6008
rect 11774 5944 11791 6008
rect 11855 5944 11872 6008
rect 11936 5944 11953 6008
rect 12017 5944 12034 6008
rect 12098 5944 12115 6008
rect 12179 5944 12196 6008
rect 12260 5944 12277 6008
rect 12341 5944 12358 6008
rect 12422 5944 12439 6008
rect 12503 5944 12520 6008
rect 12584 5944 12601 6008
rect 12665 5944 12682 6008
rect 12746 5944 12763 6008
rect 12827 5944 12844 6008
rect 12908 5944 12925 6008
rect 12989 5944 13006 6008
rect 13070 5944 13087 6008
rect 13151 5944 13168 6008
rect 13232 5944 13249 6008
rect 13313 5944 13330 6008
rect 13394 5944 13411 6008
rect 13475 5944 13492 6008
rect 13556 5944 13573 6008
rect 13637 5944 13654 6008
rect 13718 5944 13735 6008
rect 13799 5944 13816 6008
rect 13880 5944 13897 6008
rect 13961 5944 13978 6008
rect 14042 5944 14059 6008
rect 14123 5944 14140 6008
rect 14204 5944 14221 6008
rect 14285 5944 14302 6008
rect 14366 5944 14383 6008
rect 14447 5944 14464 6008
rect 14528 5944 14545 6008
rect 14609 5944 14626 6008
rect 14690 5944 14707 6008
rect 14771 5944 14788 6008
rect 14852 5944 14858 6008
rect 10078 5922 14858 5944
rect 10078 5858 10084 5922
rect 10148 5858 10166 5922
rect 10230 5858 10248 5922
rect 10312 5858 10330 5922
rect 10394 5858 10412 5922
rect 10476 5858 10494 5922
rect 10558 5858 10576 5922
rect 10640 5858 10657 5922
rect 10721 5858 10738 5922
rect 10802 5858 10819 5922
rect 10883 5858 10900 5922
rect 10964 5858 10981 5922
rect 11045 5858 11062 5922
rect 11126 5858 11143 5922
rect 11207 5858 11224 5922
rect 11288 5858 11305 5922
rect 11369 5858 11386 5922
rect 11450 5858 11467 5922
rect 11531 5858 11548 5922
rect 11612 5858 11629 5922
rect 11693 5858 11710 5922
rect 11774 5858 11791 5922
rect 11855 5858 11872 5922
rect 11936 5858 11953 5922
rect 12017 5858 12034 5922
rect 12098 5858 12115 5922
rect 12179 5858 12196 5922
rect 12260 5858 12277 5922
rect 12341 5858 12358 5922
rect 12422 5858 12439 5922
rect 12503 5858 12520 5922
rect 12584 5858 12601 5922
rect 12665 5858 12682 5922
rect 12746 5858 12763 5922
rect 12827 5858 12844 5922
rect 12908 5858 12925 5922
rect 12989 5858 13006 5922
rect 13070 5858 13087 5922
rect 13151 5858 13168 5922
rect 13232 5858 13249 5922
rect 13313 5858 13330 5922
rect 13394 5858 13411 5922
rect 13475 5858 13492 5922
rect 13556 5858 13573 5922
rect 13637 5858 13654 5922
rect 13718 5858 13735 5922
rect 13799 5858 13816 5922
rect 13880 5858 13897 5922
rect 13961 5858 13978 5922
rect 14042 5858 14059 5922
rect 14123 5858 14140 5922
rect 14204 5858 14221 5922
rect 14285 5858 14302 5922
rect 14366 5858 14383 5922
rect 14447 5858 14464 5922
rect 14528 5858 14545 5922
rect 14609 5858 14626 5922
rect 14690 5858 14707 5922
rect 14771 5858 14788 5922
rect 14852 5858 14858 5922
rect 10078 5836 14858 5858
rect 10078 5772 10084 5836
rect 10148 5772 10166 5836
rect 10230 5772 10248 5836
rect 10312 5772 10330 5836
rect 10394 5772 10412 5836
rect 10476 5772 10494 5836
rect 10558 5772 10576 5836
rect 10640 5772 10657 5836
rect 10721 5772 10738 5836
rect 10802 5772 10819 5836
rect 10883 5772 10900 5836
rect 10964 5772 10981 5836
rect 11045 5772 11062 5836
rect 11126 5772 11143 5836
rect 11207 5772 11224 5836
rect 11288 5772 11305 5836
rect 11369 5772 11386 5836
rect 11450 5772 11467 5836
rect 11531 5772 11548 5836
rect 11612 5772 11629 5836
rect 11693 5772 11710 5836
rect 11774 5772 11791 5836
rect 11855 5772 11872 5836
rect 11936 5772 11953 5836
rect 12017 5772 12034 5836
rect 12098 5772 12115 5836
rect 12179 5772 12196 5836
rect 12260 5772 12277 5836
rect 12341 5772 12358 5836
rect 12422 5772 12439 5836
rect 12503 5772 12520 5836
rect 12584 5772 12601 5836
rect 12665 5772 12682 5836
rect 12746 5772 12763 5836
rect 12827 5772 12844 5836
rect 12908 5772 12925 5836
rect 12989 5772 13006 5836
rect 13070 5772 13087 5836
rect 13151 5772 13168 5836
rect 13232 5772 13249 5836
rect 13313 5772 13330 5836
rect 13394 5772 13411 5836
rect 13475 5772 13492 5836
rect 13556 5772 13573 5836
rect 13637 5772 13654 5836
rect 13718 5772 13735 5836
rect 13799 5772 13816 5836
rect 13880 5772 13897 5836
rect 13961 5772 13978 5836
rect 14042 5772 14059 5836
rect 14123 5772 14140 5836
rect 14204 5772 14221 5836
rect 14285 5772 14302 5836
rect 14366 5772 14383 5836
rect 14447 5772 14464 5836
rect 14528 5772 14545 5836
rect 14609 5772 14626 5836
rect 14690 5772 14707 5836
rect 14771 5772 14788 5836
rect 14852 5772 14858 5836
rect 10078 5750 14858 5772
rect 10078 5686 10084 5750
rect 10148 5686 10166 5750
rect 10230 5686 10248 5750
rect 10312 5686 10330 5750
rect 10394 5686 10412 5750
rect 10476 5686 10494 5750
rect 10558 5686 10576 5750
rect 10640 5686 10657 5750
rect 10721 5686 10738 5750
rect 10802 5686 10819 5750
rect 10883 5686 10900 5750
rect 10964 5686 10981 5750
rect 11045 5686 11062 5750
rect 11126 5686 11143 5750
rect 11207 5686 11224 5750
rect 11288 5686 11305 5750
rect 11369 5686 11386 5750
rect 11450 5686 11467 5750
rect 11531 5686 11548 5750
rect 11612 5686 11629 5750
rect 11693 5686 11710 5750
rect 11774 5686 11791 5750
rect 11855 5686 11872 5750
rect 11936 5686 11953 5750
rect 12017 5686 12034 5750
rect 12098 5686 12115 5750
rect 12179 5686 12196 5750
rect 12260 5686 12277 5750
rect 12341 5686 12358 5750
rect 12422 5686 12439 5750
rect 12503 5686 12520 5750
rect 12584 5686 12601 5750
rect 12665 5686 12682 5750
rect 12746 5686 12763 5750
rect 12827 5686 12844 5750
rect 12908 5686 12925 5750
rect 12989 5686 13006 5750
rect 13070 5686 13087 5750
rect 13151 5686 13168 5750
rect 13232 5686 13249 5750
rect 13313 5686 13330 5750
rect 13394 5686 13411 5750
rect 13475 5686 13492 5750
rect 13556 5686 13573 5750
rect 13637 5686 13654 5750
rect 13718 5686 13735 5750
rect 13799 5686 13816 5750
rect 13880 5686 13897 5750
rect 13961 5686 13978 5750
rect 14042 5686 14059 5750
rect 14123 5686 14140 5750
rect 14204 5686 14221 5750
rect 14285 5686 14302 5750
rect 14366 5686 14383 5750
rect 14447 5686 14464 5750
rect 14528 5686 14545 5750
rect 14609 5686 14626 5750
rect 14690 5686 14707 5750
rect 14771 5686 14788 5750
rect 14852 5686 14858 5750
rect 10078 5664 14858 5686
rect 10078 5600 10084 5664
rect 10148 5600 10166 5664
rect 10230 5600 10248 5664
rect 10312 5600 10330 5664
rect 10394 5600 10412 5664
rect 10476 5600 10494 5664
rect 10558 5600 10576 5664
rect 10640 5600 10657 5664
rect 10721 5600 10738 5664
rect 10802 5600 10819 5664
rect 10883 5600 10900 5664
rect 10964 5600 10981 5664
rect 11045 5600 11062 5664
rect 11126 5600 11143 5664
rect 11207 5600 11224 5664
rect 11288 5600 11305 5664
rect 11369 5600 11386 5664
rect 11450 5600 11467 5664
rect 11531 5600 11548 5664
rect 11612 5600 11629 5664
rect 11693 5600 11710 5664
rect 11774 5600 11791 5664
rect 11855 5600 11872 5664
rect 11936 5600 11953 5664
rect 12017 5600 12034 5664
rect 12098 5600 12115 5664
rect 12179 5600 12196 5664
rect 12260 5600 12277 5664
rect 12341 5600 12358 5664
rect 12422 5600 12439 5664
rect 12503 5600 12520 5664
rect 12584 5600 12601 5664
rect 12665 5600 12682 5664
rect 12746 5600 12763 5664
rect 12827 5600 12844 5664
rect 12908 5600 12925 5664
rect 12989 5600 13006 5664
rect 13070 5600 13087 5664
rect 13151 5600 13168 5664
rect 13232 5600 13249 5664
rect 13313 5600 13330 5664
rect 13394 5600 13411 5664
rect 13475 5600 13492 5664
rect 13556 5600 13573 5664
rect 13637 5600 13654 5664
rect 13718 5600 13735 5664
rect 13799 5600 13816 5664
rect 13880 5600 13897 5664
rect 13961 5600 13978 5664
rect 14042 5600 14059 5664
rect 14123 5600 14140 5664
rect 14204 5600 14221 5664
rect 14285 5600 14302 5664
rect 14366 5600 14383 5664
rect 14447 5600 14464 5664
rect 14528 5600 14545 5664
rect 14609 5600 14626 5664
rect 14690 5600 14707 5664
rect 14771 5600 14788 5664
rect 14852 5600 14858 5664
rect 10078 5578 14858 5600
rect 10078 5514 10084 5578
rect 10148 5514 10166 5578
rect 10230 5514 10248 5578
rect 10312 5514 10330 5578
rect 10394 5514 10412 5578
rect 10476 5514 10494 5578
rect 10558 5514 10576 5578
rect 10640 5514 10657 5578
rect 10721 5514 10738 5578
rect 10802 5514 10819 5578
rect 10883 5514 10900 5578
rect 10964 5514 10981 5578
rect 11045 5514 11062 5578
rect 11126 5514 11143 5578
rect 11207 5514 11224 5578
rect 11288 5514 11305 5578
rect 11369 5514 11386 5578
rect 11450 5514 11467 5578
rect 11531 5514 11548 5578
rect 11612 5514 11629 5578
rect 11693 5514 11710 5578
rect 11774 5514 11791 5578
rect 11855 5514 11872 5578
rect 11936 5514 11953 5578
rect 12017 5514 12034 5578
rect 12098 5514 12115 5578
rect 12179 5514 12196 5578
rect 12260 5514 12277 5578
rect 12341 5514 12358 5578
rect 12422 5514 12439 5578
rect 12503 5514 12520 5578
rect 12584 5514 12601 5578
rect 12665 5514 12682 5578
rect 12746 5514 12763 5578
rect 12827 5514 12844 5578
rect 12908 5514 12925 5578
rect 12989 5514 13006 5578
rect 13070 5514 13087 5578
rect 13151 5514 13168 5578
rect 13232 5514 13249 5578
rect 13313 5514 13330 5578
rect 13394 5514 13411 5578
rect 13475 5514 13492 5578
rect 13556 5514 13573 5578
rect 13637 5514 13654 5578
rect 13718 5514 13735 5578
rect 13799 5514 13816 5578
rect 13880 5514 13897 5578
rect 13961 5514 13978 5578
rect 14042 5514 14059 5578
rect 14123 5514 14140 5578
rect 14204 5514 14221 5578
rect 14285 5514 14302 5578
rect 14366 5514 14383 5578
rect 14447 5514 14464 5578
rect 14528 5514 14545 5578
rect 14609 5514 14626 5578
rect 14690 5514 14707 5578
rect 14771 5514 14788 5578
rect 14852 5514 14858 5578
rect 10078 5492 14858 5514
rect 10078 5428 10084 5492
rect 10148 5428 10166 5492
rect 10230 5428 10248 5492
rect 10312 5428 10330 5492
rect 10394 5428 10412 5492
rect 10476 5428 10494 5492
rect 10558 5428 10576 5492
rect 10640 5428 10657 5492
rect 10721 5428 10738 5492
rect 10802 5428 10819 5492
rect 10883 5428 10900 5492
rect 10964 5428 10981 5492
rect 11045 5428 11062 5492
rect 11126 5428 11143 5492
rect 11207 5428 11224 5492
rect 11288 5428 11305 5492
rect 11369 5428 11386 5492
rect 11450 5428 11467 5492
rect 11531 5428 11548 5492
rect 11612 5428 11629 5492
rect 11693 5428 11710 5492
rect 11774 5428 11791 5492
rect 11855 5428 11872 5492
rect 11936 5428 11953 5492
rect 12017 5428 12034 5492
rect 12098 5428 12115 5492
rect 12179 5428 12196 5492
rect 12260 5428 12277 5492
rect 12341 5428 12358 5492
rect 12422 5428 12439 5492
rect 12503 5428 12520 5492
rect 12584 5428 12601 5492
rect 12665 5428 12682 5492
rect 12746 5428 12763 5492
rect 12827 5428 12844 5492
rect 12908 5428 12925 5492
rect 12989 5428 13006 5492
rect 13070 5428 13087 5492
rect 13151 5428 13168 5492
rect 13232 5428 13249 5492
rect 13313 5428 13330 5492
rect 13394 5428 13411 5492
rect 13475 5428 13492 5492
rect 13556 5428 13573 5492
rect 13637 5428 13654 5492
rect 13718 5428 13735 5492
rect 13799 5428 13816 5492
rect 13880 5428 13897 5492
rect 13961 5428 13978 5492
rect 14042 5428 14059 5492
rect 14123 5428 14140 5492
rect 14204 5428 14221 5492
rect 14285 5428 14302 5492
rect 14366 5428 14383 5492
rect 14447 5428 14464 5492
rect 14528 5428 14545 5492
rect 14609 5428 14626 5492
rect 14690 5428 14707 5492
rect 14771 5428 14788 5492
rect 14852 5428 14858 5492
rect 10078 5406 14858 5428
rect 10078 5342 10084 5406
rect 10148 5342 10166 5406
rect 10230 5342 10248 5406
rect 10312 5342 10330 5406
rect 10394 5342 10412 5406
rect 10476 5342 10494 5406
rect 10558 5342 10576 5406
rect 10640 5342 10657 5406
rect 10721 5342 10738 5406
rect 10802 5342 10819 5406
rect 10883 5342 10900 5406
rect 10964 5342 10981 5406
rect 11045 5342 11062 5406
rect 11126 5342 11143 5406
rect 11207 5342 11224 5406
rect 11288 5342 11305 5406
rect 11369 5342 11386 5406
rect 11450 5342 11467 5406
rect 11531 5342 11548 5406
rect 11612 5342 11629 5406
rect 11693 5342 11710 5406
rect 11774 5342 11791 5406
rect 11855 5342 11872 5406
rect 11936 5342 11953 5406
rect 12017 5342 12034 5406
rect 12098 5342 12115 5406
rect 12179 5342 12196 5406
rect 12260 5342 12277 5406
rect 12341 5342 12358 5406
rect 12422 5342 12439 5406
rect 12503 5342 12520 5406
rect 12584 5342 12601 5406
rect 12665 5342 12682 5406
rect 12746 5342 12763 5406
rect 12827 5342 12844 5406
rect 12908 5342 12925 5406
rect 12989 5342 13006 5406
rect 13070 5342 13087 5406
rect 13151 5342 13168 5406
rect 13232 5342 13249 5406
rect 13313 5342 13330 5406
rect 13394 5342 13411 5406
rect 13475 5342 13492 5406
rect 13556 5342 13573 5406
rect 13637 5342 13654 5406
rect 13718 5342 13735 5406
rect 13799 5342 13816 5406
rect 13880 5342 13897 5406
rect 13961 5342 13978 5406
rect 14042 5342 14059 5406
rect 14123 5342 14140 5406
rect 14204 5342 14221 5406
rect 14285 5342 14302 5406
rect 14366 5342 14383 5406
rect 14447 5342 14464 5406
rect 14528 5342 14545 5406
rect 14609 5342 14626 5406
rect 14690 5342 14707 5406
rect 14771 5342 14788 5406
rect 14852 5342 14858 5406
rect 10078 5320 14858 5342
rect 10078 5256 10084 5320
rect 10148 5256 10166 5320
rect 10230 5256 10248 5320
rect 10312 5256 10330 5320
rect 10394 5256 10412 5320
rect 10476 5256 10494 5320
rect 10558 5256 10576 5320
rect 10640 5256 10657 5320
rect 10721 5256 10738 5320
rect 10802 5256 10819 5320
rect 10883 5256 10900 5320
rect 10964 5256 10981 5320
rect 11045 5256 11062 5320
rect 11126 5256 11143 5320
rect 11207 5256 11224 5320
rect 11288 5256 11305 5320
rect 11369 5256 11386 5320
rect 11450 5256 11467 5320
rect 11531 5256 11548 5320
rect 11612 5256 11629 5320
rect 11693 5256 11710 5320
rect 11774 5256 11791 5320
rect 11855 5256 11872 5320
rect 11936 5256 11953 5320
rect 12017 5256 12034 5320
rect 12098 5256 12115 5320
rect 12179 5256 12196 5320
rect 12260 5256 12277 5320
rect 12341 5256 12358 5320
rect 12422 5256 12439 5320
rect 12503 5256 12520 5320
rect 12584 5256 12601 5320
rect 12665 5256 12682 5320
rect 12746 5256 12763 5320
rect 12827 5256 12844 5320
rect 12908 5256 12925 5320
rect 12989 5256 13006 5320
rect 13070 5256 13087 5320
rect 13151 5256 13168 5320
rect 13232 5256 13249 5320
rect 13313 5256 13330 5320
rect 13394 5256 13411 5320
rect 13475 5256 13492 5320
rect 13556 5256 13573 5320
rect 13637 5256 13654 5320
rect 13718 5256 13735 5320
rect 13799 5256 13816 5320
rect 13880 5256 13897 5320
rect 13961 5256 13978 5320
rect 14042 5256 14059 5320
rect 14123 5256 14140 5320
rect 14204 5256 14221 5320
rect 14285 5256 14302 5320
rect 14366 5256 14383 5320
rect 14447 5256 14464 5320
rect 14528 5256 14545 5320
rect 14609 5256 14626 5320
rect 14690 5256 14707 5320
rect 14771 5256 14788 5320
rect 14852 5256 14858 5320
rect 10078 5234 14858 5256
rect 10078 5170 10084 5234
rect 10148 5170 10166 5234
rect 10230 5170 10248 5234
rect 10312 5170 10330 5234
rect 10394 5170 10412 5234
rect 10476 5170 10494 5234
rect 10558 5170 10576 5234
rect 10640 5170 10657 5234
rect 10721 5170 10738 5234
rect 10802 5170 10819 5234
rect 10883 5170 10900 5234
rect 10964 5170 10981 5234
rect 11045 5170 11062 5234
rect 11126 5170 11143 5234
rect 11207 5170 11224 5234
rect 11288 5170 11305 5234
rect 11369 5170 11386 5234
rect 11450 5170 11467 5234
rect 11531 5170 11548 5234
rect 11612 5170 11629 5234
rect 11693 5170 11710 5234
rect 11774 5170 11791 5234
rect 11855 5170 11872 5234
rect 11936 5170 11953 5234
rect 12017 5170 12034 5234
rect 12098 5170 12115 5234
rect 12179 5170 12196 5234
rect 12260 5170 12277 5234
rect 12341 5170 12358 5234
rect 12422 5170 12439 5234
rect 12503 5170 12520 5234
rect 12584 5170 12601 5234
rect 12665 5170 12682 5234
rect 12746 5170 12763 5234
rect 12827 5170 12844 5234
rect 12908 5170 12925 5234
rect 12989 5170 13006 5234
rect 13070 5170 13087 5234
rect 13151 5170 13168 5234
rect 13232 5170 13249 5234
rect 13313 5170 13330 5234
rect 13394 5170 13411 5234
rect 13475 5170 13492 5234
rect 13556 5170 13573 5234
rect 13637 5170 13654 5234
rect 13718 5170 13735 5234
rect 13799 5170 13816 5234
rect 13880 5170 13897 5234
rect 13961 5170 13978 5234
rect 14042 5170 14059 5234
rect 14123 5170 14140 5234
rect 14204 5170 14221 5234
rect 14285 5170 14302 5234
rect 14366 5170 14383 5234
rect 14447 5170 14464 5234
rect 14528 5170 14545 5234
rect 14609 5170 14626 5234
rect 14690 5170 14707 5234
rect 14771 5170 14788 5234
rect 14852 5170 14858 5234
rect 10078 5168 14858 5170
<< via3 >>
rect 125 39919 189 39983
rect 205 39919 269 39983
rect 285 39919 349 39983
rect 365 39919 429 39983
rect 445 39919 509 39983
rect 525 39919 589 39983
rect 605 39919 669 39983
rect 685 39919 749 39983
rect 765 39919 829 39983
rect 845 39919 909 39983
rect 925 39919 989 39983
rect 1005 39919 1069 39983
rect 1085 39919 1149 39983
rect 1165 39919 1229 39983
rect 1245 39919 1309 39983
rect 1325 39919 1389 39983
rect 1405 39919 1469 39983
rect 1485 39919 1549 39983
rect 1565 39919 1629 39983
rect 1645 39919 1709 39983
rect 1725 39919 1789 39983
rect 1805 39919 1869 39983
rect 1885 39919 1949 39983
rect 1965 39919 2029 39983
rect 2045 39919 2109 39983
rect 2125 39919 2189 39983
rect 2205 39919 2269 39983
rect 2285 39919 2349 39983
rect 2365 39919 2429 39983
rect 2445 39919 2509 39983
rect 2525 39919 2589 39983
rect 2605 39919 2669 39983
rect 2727 39918 2791 39982
rect 2808 39918 2872 39982
rect 2889 39918 2953 39982
rect 2970 39918 3034 39982
rect 3051 39918 3115 39982
rect 3132 39918 3196 39982
rect 3213 39918 3277 39982
rect 3294 39918 3358 39982
rect 3375 39918 3439 39982
rect 3456 39918 3520 39982
rect 3537 39918 3601 39982
rect 3618 39918 3682 39982
rect 3699 39918 3763 39982
rect 3780 39918 3844 39982
rect 3861 39918 3925 39982
rect 3942 39918 4006 39982
rect 4023 39918 4087 39982
rect 4104 39918 4168 39982
rect 4185 39918 4249 39982
rect 4266 39918 4330 39982
rect 4347 39918 4411 39982
rect 4428 39918 4492 39982
rect 4509 39918 4573 39982
rect 4590 39918 4654 39982
rect 4671 39918 4735 39982
rect 4752 39918 4816 39982
rect 4833 39918 4897 39982
rect 4914 39918 4978 39982
rect 4995 39918 5059 39982
rect 5076 39918 5140 39982
rect 5157 39918 5221 39982
rect 5238 39918 5302 39982
rect 5319 39918 5383 39982
rect 125 39838 189 39902
rect 205 39838 269 39902
rect 285 39838 349 39902
rect 365 39838 429 39902
rect 445 39838 509 39902
rect 525 39838 589 39902
rect 605 39838 669 39902
rect 685 39838 749 39902
rect 765 39838 829 39902
rect 845 39838 909 39902
rect 925 39838 989 39902
rect 1005 39838 1069 39902
rect 1085 39838 1149 39902
rect 1165 39838 1229 39902
rect 1245 39838 1309 39902
rect 1325 39838 1389 39902
rect 1405 39838 1469 39902
rect 1485 39838 1549 39902
rect 1565 39838 1629 39902
rect 1645 39838 1709 39902
rect 1725 39838 1789 39902
rect 1805 39838 1869 39902
rect 1885 39838 1949 39902
rect 1965 39838 2029 39902
rect 2045 39838 2109 39902
rect 2125 39838 2189 39902
rect 2205 39838 2269 39902
rect 2285 39838 2349 39902
rect 2365 39838 2429 39902
rect 2445 39838 2509 39902
rect 2525 39838 2589 39902
rect 2605 39838 2669 39902
rect 2727 39838 2791 39902
rect 2808 39838 2872 39902
rect 2889 39838 2953 39902
rect 2970 39838 3034 39902
rect 3051 39838 3115 39902
rect 3132 39838 3196 39902
rect 3213 39838 3277 39902
rect 3294 39838 3358 39902
rect 3375 39838 3439 39902
rect 3456 39838 3520 39902
rect 3537 39838 3601 39902
rect 3618 39838 3682 39902
rect 3699 39838 3763 39902
rect 3780 39838 3844 39902
rect 3861 39838 3925 39902
rect 3942 39838 4006 39902
rect 4023 39838 4087 39902
rect 4104 39838 4168 39902
rect 4185 39838 4249 39902
rect 4266 39838 4330 39902
rect 4347 39838 4411 39902
rect 4428 39838 4492 39902
rect 4509 39838 4573 39902
rect 4590 39838 4654 39902
rect 4671 39838 4735 39902
rect 4752 39838 4816 39902
rect 4833 39838 4897 39902
rect 4914 39838 4978 39902
rect 4995 39838 5059 39902
rect 5076 39838 5140 39902
rect 5157 39838 5221 39902
rect 5238 39838 5302 39902
rect 5319 39838 5383 39902
rect 125 39757 189 39821
rect 205 39757 269 39821
rect 285 39757 349 39821
rect 365 39757 429 39821
rect 445 39757 509 39821
rect 525 39757 589 39821
rect 605 39757 669 39821
rect 685 39757 749 39821
rect 765 39757 829 39821
rect 845 39757 909 39821
rect 925 39757 989 39821
rect 1005 39757 1069 39821
rect 1085 39757 1149 39821
rect 1165 39757 1229 39821
rect 1245 39757 1309 39821
rect 1325 39757 1389 39821
rect 1405 39757 1469 39821
rect 1485 39757 1549 39821
rect 1565 39757 1629 39821
rect 1645 39757 1709 39821
rect 1725 39757 1789 39821
rect 1805 39757 1869 39821
rect 1885 39757 1949 39821
rect 1965 39757 2029 39821
rect 2045 39757 2109 39821
rect 2125 39757 2189 39821
rect 2205 39757 2269 39821
rect 2285 39757 2349 39821
rect 2365 39757 2429 39821
rect 2445 39757 2509 39821
rect 2525 39757 2589 39821
rect 2605 39757 2669 39821
rect 2727 39758 2791 39822
rect 2808 39758 2872 39822
rect 2889 39758 2953 39822
rect 2970 39758 3034 39822
rect 3051 39758 3115 39822
rect 3132 39758 3196 39822
rect 3213 39758 3277 39822
rect 3294 39758 3358 39822
rect 3375 39758 3439 39822
rect 3456 39758 3520 39822
rect 3537 39758 3601 39822
rect 3618 39758 3682 39822
rect 3699 39758 3763 39822
rect 3780 39758 3844 39822
rect 3861 39758 3925 39822
rect 3942 39758 4006 39822
rect 4023 39758 4087 39822
rect 4104 39758 4168 39822
rect 4185 39758 4249 39822
rect 4266 39758 4330 39822
rect 4347 39758 4411 39822
rect 4428 39758 4492 39822
rect 4509 39758 4573 39822
rect 4590 39758 4654 39822
rect 4671 39758 4735 39822
rect 4752 39758 4816 39822
rect 4833 39758 4897 39822
rect 4914 39758 4978 39822
rect 4995 39758 5059 39822
rect 5076 39758 5140 39822
rect 5157 39758 5221 39822
rect 5238 39758 5302 39822
rect 5319 39758 5383 39822
rect 125 39676 189 39740
rect 205 39676 269 39740
rect 285 39676 349 39740
rect 365 39676 429 39740
rect 445 39676 509 39740
rect 525 39676 589 39740
rect 605 39676 669 39740
rect 685 39676 749 39740
rect 765 39676 829 39740
rect 845 39676 909 39740
rect 925 39676 989 39740
rect 1005 39676 1069 39740
rect 1085 39676 1149 39740
rect 1165 39676 1229 39740
rect 1245 39676 1309 39740
rect 1325 39676 1389 39740
rect 1405 39676 1469 39740
rect 1485 39676 1549 39740
rect 1565 39676 1629 39740
rect 1645 39676 1709 39740
rect 1725 39676 1789 39740
rect 1805 39676 1869 39740
rect 1885 39676 1949 39740
rect 1965 39676 2029 39740
rect 2045 39676 2109 39740
rect 2125 39676 2189 39740
rect 2205 39676 2269 39740
rect 2285 39676 2349 39740
rect 2365 39676 2429 39740
rect 2445 39676 2509 39740
rect 2525 39676 2589 39740
rect 2605 39676 2669 39740
rect 2727 39678 2791 39742
rect 2808 39678 2872 39742
rect 2889 39678 2953 39742
rect 2970 39678 3034 39742
rect 3051 39678 3115 39742
rect 3132 39678 3196 39742
rect 3213 39678 3277 39742
rect 3294 39678 3358 39742
rect 3375 39678 3439 39742
rect 3456 39678 3520 39742
rect 3537 39678 3601 39742
rect 3618 39678 3682 39742
rect 3699 39678 3763 39742
rect 3780 39678 3844 39742
rect 3861 39678 3925 39742
rect 3942 39678 4006 39742
rect 4023 39678 4087 39742
rect 4104 39678 4168 39742
rect 4185 39678 4249 39742
rect 4266 39678 4330 39742
rect 4347 39678 4411 39742
rect 4428 39678 4492 39742
rect 4509 39678 4573 39742
rect 4590 39678 4654 39742
rect 4671 39678 4735 39742
rect 4752 39678 4816 39742
rect 4833 39678 4897 39742
rect 4914 39678 4978 39742
rect 4995 39678 5059 39742
rect 5076 39678 5140 39742
rect 5157 39678 5221 39742
rect 5238 39678 5302 39742
rect 5319 39678 5383 39742
rect 125 39595 189 39659
rect 205 39595 269 39659
rect 285 39595 349 39659
rect 365 39595 429 39659
rect 445 39595 509 39659
rect 525 39595 589 39659
rect 605 39595 669 39659
rect 685 39595 749 39659
rect 765 39595 829 39659
rect 845 39595 909 39659
rect 925 39595 989 39659
rect 1005 39595 1069 39659
rect 1085 39595 1149 39659
rect 1165 39595 1229 39659
rect 1245 39595 1309 39659
rect 1325 39595 1389 39659
rect 1405 39595 1469 39659
rect 1485 39595 1549 39659
rect 1565 39595 1629 39659
rect 1645 39595 1709 39659
rect 1725 39595 1789 39659
rect 1805 39595 1869 39659
rect 1885 39595 1949 39659
rect 1965 39595 2029 39659
rect 2045 39595 2109 39659
rect 2125 39595 2189 39659
rect 2205 39595 2269 39659
rect 2285 39595 2349 39659
rect 2365 39595 2429 39659
rect 2445 39595 2509 39659
rect 2525 39595 2589 39659
rect 2605 39595 2669 39659
rect 2727 39598 2791 39662
rect 2808 39598 2872 39662
rect 2889 39598 2953 39662
rect 2970 39598 3034 39662
rect 3051 39598 3115 39662
rect 3132 39598 3196 39662
rect 3213 39598 3277 39662
rect 3294 39598 3358 39662
rect 3375 39598 3439 39662
rect 3456 39598 3520 39662
rect 3537 39598 3601 39662
rect 3618 39598 3682 39662
rect 3699 39598 3763 39662
rect 3780 39598 3844 39662
rect 3861 39598 3925 39662
rect 3942 39598 4006 39662
rect 4023 39598 4087 39662
rect 4104 39598 4168 39662
rect 4185 39598 4249 39662
rect 4266 39598 4330 39662
rect 4347 39598 4411 39662
rect 4428 39598 4492 39662
rect 4509 39598 4573 39662
rect 4590 39598 4654 39662
rect 4671 39598 4735 39662
rect 4752 39598 4816 39662
rect 4833 39598 4897 39662
rect 4914 39598 4978 39662
rect 4995 39598 5059 39662
rect 5076 39598 5140 39662
rect 5157 39598 5221 39662
rect 5238 39598 5302 39662
rect 5319 39598 5383 39662
rect 125 39514 189 39578
rect 205 39514 269 39578
rect 285 39514 349 39578
rect 365 39514 429 39578
rect 445 39514 509 39578
rect 525 39514 589 39578
rect 605 39514 669 39578
rect 685 39514 749 39578
rect 765 39514 829 39578
rect 845 39514 909 39578
rect 925 39514 989 39578
rect 1005 39514 1069 39578
rect 1085 39514 1149 39578
rect 1165 39514 1229 39578
rect 1245 39514 1309 39578
rect 1325 39514 1389 39578
rect 1405 39514 1469 39578
rect 1485 39514 1549 39578
rect 1565 39514 1629 39578
rect 1645 39514 1709 39578
rect 1725 39514 1789 39578
rect 1805 39514 1869 39578
rect 1885 39514 1949 39578
rect 1965 39514 2029 39578
rect 2045 39514 2109 39578
rect 2125 39514 2189 39578
rect 2205 39514 2269 39578
rect 2285 39514 2349 39578
rect 2365 39514 2429 39578
rect 2445 39514 2509 39578
rect 2525 39514 2589 39578
rect 2605 39514 2669 39578
rect 2727 39518 2791 39582
rect 2808 39518 2872 39582
rect 2889 39518 2953 39582
rect 2970 39518 3034 39582
rect 3051 39518 3115 39582
rect 3132 39518 3196 39582
rect 3213 39518 3277 39582
rect 3294 39518 3358 39582
rect 3375 39518 3439 39582
rect 3456 39518 3520 39582
rect 3537 39518 3601 39582
rect 3618 39518 3682 39582
rect 3699 39518 3763 39582
rect 3780 39518 3844 39582
rect 3861 39518 3925 39582
rect 3942 39518 4006 39582
rect 4023 39518 4087 39582
rect 4104 39518 4168 39582
rect 4185 39518 4249 39582
rect 4266 39518 4330 39582
rect 4347 39518 4411 39582
rect 4428 39518 4492 39582
rect 4509 39518 4573 39582
rect 4590 39518 4654 39582
rect 4671 39518 4735 39582
rect 4752 39518 4816 39582
rect 4833 39518 4897 39582
rect 4914 39518 4978 39582
rect 4995 39518 5059 39582
rect 5076 39518 5140 39582
rect 5157 39518 5221 39582
rect 5238 39518 5302 39582
rect 5319 39518 5383 39582
rect 125 39433 189 39497
rect 205 39433 269 39497
rect 285 39433 349 39497
rect 365 39433 429 39497
rect 445 39433 509 39497
rect 525 39433 589 39497
rect 605 39433 669 39497
rect 685 39433 749 39497
rect 765 39433 829 39497
rect 845 39433 909 39497
rect 925 39433 989 39497
rect 1005 39433 1069 39497
rect 1085 39433 1149 39497
rect 1165 39433 1229 39497
rect 1245 39433 1309 39497
rect 1325 39433 1389 39497
rect 1405 39433 1469 39497
rect 1485 39433 1549 39497
rect 1565 39433 1629 39497
rect 1645 39433 1709 39497
rect 1725 39433 1789 39497
rect 1805 39433 1869 39497
rect 1885 39433 1949 39497
rect 1965 39433 2029 39497
rect 2045 39433 2109 39497
rect 2125 39433 2189 39497
rect 2205 39433 2269 39497
rect 2285 39433 2349 39497
rect 2365 39433 2429 39497
rect 2445 39433 2509 39497
rect 2525 39433 2589 39497
rect 2605 39433 2669 39497
rect 2727 39438 2791 39502
rect 2808 39438 2872 39502
rect 2889 39438 2953 39502
rect 2970 39438 3034 39502
rect 3051 39438 3115 39502
rect 3132 39438 3196 39502
rect 3213 39438 3277 39502
rect 3294 39438 3358 39502
rect 3375 39438 3439 39502
rect 3456 39438 3520 39502
rect 3537 39438 3601 39502
rect 3618 39438 3682 39502
rect 3699 39438 3763 39502
rect 3780 39438 3844 39502
rect 3861 39438 3925 39502
rect 3942 39438 4006 39502
rect 4023 39438 4087 39502
rect 4104 39438 4168 39502
rect 4185 39438 4249 39502
rect 4266 39438 4330 39502
rect 4347 39438 4411 39502
rect 4428 39438 4492 39502
rect 4509 39438 4573 39502
rect 4590 39438 4654 39502
rect 4671 39438 4735 39502
rect 4752 39438 4816 39502
rect 4833 39438 4897 39502
rect 4914 39438 4978 39502
rect 4995 39438 5059 39502
rect 5076 39438 5140 39502
rect 5157 39438 5221 39502
rect 5238 39438 5302 39502
rect 5319 39438 5383 39502
rect 5400 39438 12264 39982
rect 12306 39919 12370 39983
rect 12386 39919 12450 39983
rect 12466 39919 12530 39983
rect 12546 39919 12610 39983
rect 12626 39919 12690 39983
rect 12706 39919 12770 39983
rect 12786 39919 12850 39983
rect 12866 39919 12930 39983
rect 12946 39919 13010 39983
rect 13026 39919 13090 39983
rect 13106 39919 13170 39983
rect 13186 39919 13250 39983
rect 13266 39919 13330 39983
rect 13346 39919 13410 39983
rect 13426 39919 13490 39983
rect 13506 39919 13570 39983
rect 13586 39919 13650 39983
rect 13666 39919 13730 39983
rect 13746 39919 13810 39983
rect 13826 39919 13890 39983
rect 13906 39919 13970 39983
rect 13986 39919 14050 39983
rect 14066 39919 14130 39983
rect 14146 39919 14210 39983
rect 14226 39919 14290 39983
rect 14306 39919 14370 39983
rect 14386 39919 14450 39983
rect 14466 39919 14530 39983
rect 14546 39919 14610 39983
rect 14626 39919 14690 39983
rect 14706 39919 14770 39983
rect 14786 39919 14850 39983
rect 12306 39838 12370 39902
rect 12386 39838 12450 39902
rect 12466 39838 12530 39902
rect 12546 39838 12610 39902
rect 12626 39838 12690 39902
rect 12706 39838 12770 39902
rect 12786 39838 12850 39902
rect 12866 39838 12930 39902
rect 12946 39838 13010 39902
rect 13026 39838 13090 39902
rect 13106 39838 13170 39902
rect 13186 39838 13250 39902
rect 13266 39838 13330 39902
rect 13346 39838 13410 39902
rect 13426 39838 13490 39902
rect 13506 39838 13570 39902
rect 13586 39838 13650 39902
rect 13666 39838 13730 39902
rect 13746 39838 13810 39902
rect 13826 39838 13890 39902
rect 13906 39838 13970 39902
rect 13986 39838 14050 39902
rect 14066 39838 14130 39902
rect 14146 39838 14210 39902
rect 14226 39838 14290 39902
rect 14306 39838 14370 39902
rect 14386 39838 14450 39902
rect 14466 39838 14530 39902
rect 14546 39838 14610 39902
rect 14626 39838 14690 39902
rect 14706 39838 14770 39902
rect 14786 39838 14850 39902
rect 12306 39757 12370 39821
rect 12386 39757 12450 39821
rect 12466 39757 12530 39821
rect 12546 39757 12610 39821
rect 12626 39757 12690 39821
rect 12706 39757 12770 39821
rect 12786 39757 12850 39821
rect 12866 39757 12930 39821
rect 12946 39757 13010 39821
rect 13026 39757 13090 39821
rect 13106 39757 13170 39821
rect 13186 39757 13250 39821
rect 13266 39757 13330 39821
rect 13346 39757 13410 39821
rect 13426 39757 13490 39821
rect 13506 39757 13570 39821
rect 13586 39757 13650 39821
rect 13666 39757 13730 39821
rect 13746 39757 13810 39821
rect 13826 39757 13890 39821
rect 13906 39757 13970 39821
rect 13986 39757 14050 39821
rect 14066 39757 14130 39821
rect 14146 39757 14210 39821
rect 14226 39757 14290 39821
rect 14306 39757 14370 39821
rect 14386 39757 14450 39821
rect 14466 39757 14530 39821
rect 14546 39757 14610 39821
rect 14626 39757 14690 39821
rect 14706 39757 14770 39821
rect 14786 39757 14850 39821
rect 12306 39676 12370 39740
rect 12386 39676 12450 39740
rect 12466 39676 12530 39740
rect 12546 39676 12610 39740
rect 12626 39676 12690 39740
rect 12706 39676 12770 39740
rect 12786 39676 12850 39740
rect 12866 39676 12930 39740
rect 12946 39676 13010 39740
rect 13026 39676 13090 39740
rect 13106 39676 13170 39740
rect 13186 39676 13250 39740
rect 13266 39676 13330 39740
rect 13346 39676 13410 39740
rect 13426 39676 13490 39740
rect 13506 39676 13570 39740
rect 13586 39676 13650 39740
rect 13666 39676 13730 39740
rect 13746 39676 13810 39740
rect 13826 39676 13890 39740
rect 13906 39676 13970 39740
rect 13986 39676 14050 39740
rect 14066 39676 14130 39740
rect 14146 39676 14210 39740
rect 14226 39676 14290 39740
rect 14306 39676 14370 39740
rect 14386 39676 14450 39740
rect 14466 39676 14530 39740
rect 14546 39676 14610 39740
rect 14626 39676 14690 39740
rect 14706 39676 14770 39740
rect 14786 39676 14850 39740
rect 12306 39595 12370 39659
rect 12386 39595 12450 39659
rect 12466 39595 12530 39659
rect 12546 39595 12610 39659
rect 12626 39595 12690 39659
rect 12706 39595 12770 39659
rect 12786 39595 12850 39659
rect 12866 39595 12930 39659
rect 12946 39595 13010 39659
rect 13026 39595 13090 39659
rect 13106 39595 13170 39659
rect 13186 39595 13250 39659
rect 13266 39595 13330 39659
rect 13346 39595 13410 39659
rect 13426 39595 13490 39659
rect 13506 39595 13570 39659
rect 13586 39595 13650 39659
rect 13666 39595 13730 39659
rect 13746 39595 13810 39659
rect 13826 39595 13890 39659
rect 13906 39595 13970 39659
rect 13986 39595 14050 39659
rect 14066 39595 14130 39659
rect 14146 39595 14210 39659
rect 14226 39595 14290 39659
rect 14306 39595 14370 39659
rect 14386 39595 14450 39659
rect 14466 39595 14530 39659
rect 14546 39595 14610 39659
rect 14626 39595 14690 39659
rect 14706 39595 14770 39659
rect 14786 39595 14850 39659
rect 12306 39514 12370 39578
rect 12386 39514 12450 39578
rect 12466 39514 12530 39578
rect 12546 39514 12610 39578
rect 12626 39514 12690 39578
rect 12706 39514 12770 39578
rect 12786 39514 12850 39578
rect 12866 39514 12930 39578
rect 12946 39514 13010 39578
rect 13026 39514 13090 39578
rect 13106 39514 13170 39578
rect 13186 39514 13250 39578
rect 13266 39514 13330 39578
rect 13346 39514 13410 39578
rect 13426 39514 13490 39578
rect 13506 39514 13570 39578
rect 13586 39514 13650 39578
rect 13666 39514 13730 39578
rect 13746 39514 13810 39578
rect 13826 39514 13890 39578
rect 13906 39514 13970 39578
rect 13986 39514 14050 39578
rect 14066 39514 14130 39578
rect 14146 39514 14210 39578
rect 14226 39514 14290 39578
rect 14306 39514 14370 39578
rect 14386 39514 14450 39578
rect 14466 39514 14530 39578
rect 14546 39514 14610 39578
rect 14626 39514 14690 39578
rect 14706 39514 14770 39578
rect 14786 39514 14850 39578
rect 125 39352 189 39416
rect 205 39352 269 39416
rect 285 39352 349 39416
rect 365 39352 429 39416
rect 445 39352 509 39416
rect 525 39352 589 39416
rect 605 39352 669 39416
rect 685 39352 749 39416
rect 765 39352 829 39416
rect 845 39352 909 39416
rect 925 39352 989 39416
rect 1005 39352 1069 39416
rect 1085 39352 1149 39416
rect 1165 39352 1229 39416
rect 1245 39352 1309 39416
rect 1325 39352 1389 39416
rect 1405 39352 1469 39416
rect 1485 39352 1549 39416
rect 1565 39352 1629 39416
rect 1645 39352 1709 39416
rect 1725 39352 1789 39416
rect 1805 39352 1869 39416
rect 1885 39352 1949 39416
rect 1965 39352 2029 39416
rect 2045 39352 2109 39416
rect 2125 39352 2189 39416
rect 2205 39352 2269 39416
rect 2285 39352 2349 39416
rect 2365 39352 2429 39416
rect 2445 39352 2509 39416
rect 2525 39352 2589 39416
rect 2605 39352 2669 39416
rect 12306 39433 12370 39497
rect 12386 39433 12450 39497
rect 12466 39433 12530 39497
rect 12546 39433 12610 39497
rect 12626 39433 12690 39497
rect 12706 39433 12770 39497
rect 12786 39433 12850 39497
rect 12866 39433 12930 39497
rect 12946 39433 13010 39497
rect 13026 39433 13090 39497
rect 13106 39433 13170 39497
rect 13186 39433 13250 39497
rect 13266 39433 13330 39497
rect 13346 39433 13410 39497
rect 13426 39433 13490 39497
rect 13506 39433 13570 39497
rect 13586 39433 13650 39497
rect 13666 39433 13730 39497
rect 13746 39433 13810 39497
rect 13826 39433 13890 39497
rect 13906 39433 13970 39497
rect 13986 39433 14050 39497
rect 14066 39433 14130 39497
rect 14146 39433 14210 39497
rect 14226 39433 14290 39497
rect 14306 39433 14370 39497
rect 14386 39433 14450 39497
rect 14466 39433 14530 39497
rect 14546 39433 14610 39497
rect 14626 39433 14690 39497
rect 14706 39433 14770 39497
rect 14786 39433 14850 39497
rect 125 39271 189 39335
rect 205 39271 269 39335
rect 285 39271 349 39335
rect 365 39271 429 39335
rect 445 39271 509 39335
rect 525 39271 589 39335
rect 605 39271 669 39335
rect 685 39271 749 39335
rect 765 39271 829 39335
rect 845 39271 909 39335
rect 925 39271 989 39335
rect 1005 39271 1069 39335
rect 1085 39271 1149 39335
rect 1165 39271 1229 39335
rect 1245 39271 1309 39335
rect 1325 39271 1389 39335
rect 1405 39271 1469 39335
rect 1485 39271 1549 39335
rect 1565 39271 1629 39335
rect 1645 39271 1709 39335
rect 1725 39271 1789 39335
rect 1805 39271 1869 39335
rect 1885 39271 1949 39335
rect 1965 39271 2029 39335
rect 2045 39271 2109 39335
rect 2125 39271 2189 39335
rect 2205 39271 2269 39335
rect 2285 39271 2349 39335
rect 2365 39271 2429 39335
rect 2445 39271 2509 39335
rect 2525 39271 2589 39335
rect 2605 39271 2669 39335
rect 2753 39329 2817 39393
rect 125 39190 189 39254
rect 205 39190 269 39254
rect 285 39190 349 39254
rect 365 39190 429 39254
rect 445 39190 509 39254
rect 525 39190 589 39254
rect 605 39190 669 39254
rect 685 39190 749 39254
rect 765 39190 829 39254
rect 845 39190 909 39254
rect 925 39190 989 39254
rect 1005 39190 1069 39254
rect 1085 39190 1149 39254
rect 1165 39190 1229 39254
rect 1245 39190 1309 39254
rect 1325 39190 1389 39254
rect 1405 39190 1469 39254
rect 1485 39190 1549 39254
rect 1565 39190 1629 39254
rect 1645 39190 1709 39254
rect 1725 39190 1789 39254
rect 1805 39190 1869 39254
rect 1885 39190 1949 39254
rect 1965 39190 2029 39254
rect 2045 39190 2109 39254
rect 2125 39190 2189 39254
rect 2205 39190 2269 39254
rect 2285 39190 2349 39254
rect 2365 39190 2429 39254
rect 2445 39190 2509 39254
rect 2525 39190 2589 39254
rect 2605 39190 2669 39254
rect 2753 39247 2817 39311
rect 12170 39329 12234 39393
rect 12306 39352 12370 39416
rect 12386 39352 12450 39416
rect 12466 39352 12530 39416
rect 12546 39352 12610 39416
rect 12626 39352 12690 39416
rect 12706 39352 12770 39416
rect 12786 39352 12850 39416
rect 12866 39352 12930 39416
rect 12946 39352 13010 39416
rect 13026 39352 13090 39416
rect 13106 39352 13170 39416
rect 13186 39352 13250 39416
rect 13266 39352 13330 39416
rect 13346 39352 13410 39416
rect 13426 39352 13490 39416
rect 13506 39352 13570 39416
rect 13586 39352 13650 39416
rect 13666 39352 13730 39416
rect 13746 39352 13810 39416
rect 13826 39352 13890 39416
rect 13906 39352 13970 39416
rect 13986 39352 14050 39416
rect 14066 39352 14130 39416
rect 14146 39352 14210 39416
rect 14226 39352 14290 39416
rect 14306 39352 14370 39416
rect 14386 39352 14450 39416
rect 14466 39352 14530 39416
rect 14546 39352 14610 39416
rect 14626 39352 14690 39416
rect 14706 39352 14770 39416
rect 14786 39352 14850 39416
rect 12170 39247 12234 39311
rect 12306 39271 12370 39335
rect 12386 39271 12450 39335
rect 12466 39271 12530 39335
rect 12546 39271 12610 39335
rect 12626 39271 12690 39335
rect 12706 39271 12770 39335
rect 12786 39271 12850 39335
rect 12866 39271 12930 39335
rect 12946 39271 13010 39335
rect 13026 39271 13090 39335
rect 13106 39271 13170 39335
rect 13186 39271 13250 39335
rect 13266 39271 13330 39335
rect 13346 39271 13410 39335
rect 13426 39271 13490 39335
rect 13506 39271 13570 39335
rect 13586 39271 13650 39335
rect 13666 39271 13730 39335
rect 13746 39271 13810 39335
rect 13826 39271 13890 39335
rect 13906 39271 13970 39335
rect 13986 39271 14050 39335
rect 14066 39271 14130 39335
rect 14146 39271 14210 39335
rect 14226 39271 14290 39335
rect 14306 39271 14370 39335
rect 14386 39271 14450 39335
rect 14466 39271 14530 39335
rect 14546 39271 14610 39335
rect 14626 39271 14690 39335
rect 14706 39271 14770 39335
rect 14786 39271 14850 39335
rect 125 39109 189 39173
rect 205 39109 269 39173
rect 285 39109 349 39173
rect 365 39109 429 39173
rect 445 39109 509 39173
rect 525 39109 589 39173
rect 605 39109 669 39173
rect 685 39109 749 39173
rect 765 39109 829 39173
rect 845 39109 909 39173
rect 925 39109 989 39173
rect 1005 39109 1069 39173
rect 1085 39109 1149 39173
rect 1165 39109 1229 39173
rect 1245 39109 1309 39173
rect 1325 39109 1389 39173
rect 1405 39109 1469 39173
rect 1485 39109 1549 39173
rect 1565 39109 1629 39173
rect 1645 39109 1709 39173
rect 1725 39109 1789 39173
rect 1805 39109 1869 39173
rect 1885 39109 1949 39173
rect 1965 39109 2029 39173
rect 2045 39109 2109 39173
rect 2125 39109 2189 39173
rect 2205 39109 2269 39173
rect 2285 39109 2349 39173
rect 2365 39109 2429 39173
rect 2445 39109 2509 39173
rect 2525 39109 2589 39173
rect 2605 39109 2669 39173
rect 125 39028 189 39092
rect 205 39028 269 39092
rect 285 39028 349 39092
rect 365 39028 429 39092
rect 445 39028 509 39092
rect 525 39028 589 39092
rect 605 39028 669 39092
rect 685 39028 749 39092
rect 765 39028 829 39092
rect 845 39028 909 39092
rect 925 39028 989 39092
rect 1005 39028 1069 39092
rect 1085 39028 1149 39092
rect 1165 39028 1229 39092
rect 1245 39028 1309 39092
rect 1325 39028 1389 39092
rect 1405 39028 1469 39092
rect 1485 39028 1549 39092
rect 1565 39028 1629 39092
rect 1645 39028 1709 39092
rect 1725 39028 1789 39092
rect 1805 39028 1869 39092
rect 1885 39028 1949 39092
rect 1965 39028 2029 39092
rect 2045 39028 2109 39092
rect 2125 39028 2189 39092
rect 2205 39028 2269 39092
rect 2285 39028 2349 39092
rect 2365 39028 2429 39092
rect 2445 39028 2509 39092
rect 2525 39028 2589 39092
rect 2605 39028 2669 39092
rect 12306 39190 12370 39254
rect 12386 39190 12450 39254
rect 12466 39190 12530 39254
rect 12546 39190 12610 39254
rect 12626 39190 12690 39254
rect 12706 39190 12770 39254
rect 12786 39190 12850 39254
rect 12866 39190 12930 39254
rect 12946 39190 13010 39254
rect 13026 39190 13090 39254
rect 13106 39190 13170 39254
rect 13186 39190 13250 39254
rect 13266 39190 13330 39254
rect 13346 39190 13410 39254
rect 13426 39190 13490 39254
rect 13506 39190 13570 39254
rect 13586 39190 13650 39254
rect 13666 39190 13730 39254
rect 13746 39190 13810 39254
rect 13826 39190 13890 39254
rect 13906 39190 13970 39254
rect 13986 39190 14050 39254
rect 14066 39190 14130 39254
rect 14146 39190 14210 39254
rect 14226 39190 14290 39254
rect 14306 39190 14370 39254
rect 14386 39190 14450 39254
rect 14466 39190 14530 39254
rect 14546 39190 14610 39254
rect 14626 39190 14690 39254
rect 14706 39190 14770 39254
rect 14786 39190 14850 39254
rect 12306 39109 12370 39173
rect 12386 39109 12450 39173
rect 12466 39109 12530 39173
rect 12546 39109 12610 39173
rect 12626 39109 12690 39173
rect 12706 39109 12770 39173
rect 12786 39109 12850 39173
rect 12866 39109 12930 39173
rect 12946 39109 13010 39173
rect 13026 39109 13090 39173
rect 13106 39109 13170 39173
rect 13186 39109 13250 39173
rect 13266 39109 13330 39173
rect 13346 39109 13410 39173
rect 13426 39109 13490 39173
rect 13506 39109 13570 39173
rect 13586 39109 13650 39173
rect 13666 39109 13730 39173
rect 13746 39109 13810 39173
rect 13826 39109 13890 39173
rect 13906 39109 13970 39173
rect 13986 39109 14050 39173
rect 14066 39109 14130 39173
rect 14146 39109 14210 39173
rect 14226 39109 14290 39173
rect 14306 39109 14370 39173
rect 14386 39109 14450 39173
rect 14466 39109 14530 39173
rect 14546 39109 14610 39173
rect 14626 39109 14690 39173
rect 14706 39109 14770 39173
rect 14786 39109 14850 39173
rect 125 35187 2669 39011
rect 12306 39028 12370 39092
rect 12386 39028 12450 39092
rect 12466 39028 12530 39092
rect 12546 39028 12610 39092
rect 12626 39028 12690 39092
rect 12706 39028 12770 39092
rect 12786 39028 12850 39092
rect 12866 39028 12930 39092
rect 12946 39028 13010 39092
rect 13026 39028 13090 39092
rect 13106 39028 13170 39092
rect 13186 39028 13250 39092
rect 13266 39028 13330 39092
rect 13346 39028 13410 39092
rect 13426 39028 13490 39092
rect 13506 39028 13570 39092
rect 13586 39028 13650 39092
rect 13666 39028 13730 39092
rect 13746 39028 13810 39092
rect 13826 39028 13890 39092
rect 13906 39028 13970 39092
rect 13986 39028 14050 39092
rect 14066 39028 14130 39092
rect 14146 39028 14210 39092
rect 14226 39028 14290 39092
rect 14306 39028 14370 39092
rect 14386 39028 14450 39092
rect 14466 39028 14530 39092
rect 14546 39028 14610 39092
rect 14626 39028 14690 39092
rect 14706 39028 14770 39092
rect 14786 39028 14850 39092
rect 12306 35187 14850 39011
rect 105 12470 169 12534
rect 187 12470 251 12534
rect 269 12470 333 12534
rect 351 12470 415 12534
rect 433 12470 497 12534
rect 515 12470 579 12534
rect 597 12470 661 12534
rect 678 12470 742 12534
rect 759 12470 823 12534
rect 840 12470 904 12534
rect 921 12470 985 12534
rect 1002 12470 1066 12534
rect 1083 12470 1147 12534
rect 1164 12470 1228 12534
rect 1245 12470 1309 12534
rect 1326 12470 1390 12534
rect 1407 12470 1471 12534
rect 1488 12470 1552 12534
rect 1569 12470 1633 12534
rect 1650 12470 1714 12534
rect 1731 12470 1795 12534
rect 1812 12470 1876 12534
rect 1893 12470 1957 12534
rect 1974 12470 2038 12534
rect 2055 12470 2119 12534
rect 2136 12470 2200 12534
rect 2217 12470 2281 12534
rect 2298 12470 2362 12534
rect 2379 12470 2443 12534
rect 2460 12470 2524 12534
rect 2541 12470 2605 12534
rect 2622 12470 2686 12534
rect 2703 12470 2767 12534
rect 2784 12470 2848 12534
rect 2865 12470 2929 12534
rect 2946 12470 3010 12534
rect 3027 12470 3091 12534
rect 3108 12470 3172 12534
rect 3189 12470 3253 12534
rect 3270 12470 3334 12534
rect 3351 12470 3415 12534
rect 3432 12470 3496 12534
rect 3513 12470 3577 12534
rect 3594 12470 3658 12534
rect 3675 12470 3739 12534
rect 3756 12470 3820 12534
rect 3837 12470 3901 12534
rect 3918 12470 3982 12534
rect 3999 12470 4063 12534
rect 4080 12470 4144 12534
rect 4161 12470 4225 12534
rect 4242 12470 4306 12534
rect 4323 12470 4387 12534
rect 4404 12470 4468 12534
rect 4485 12470 4549 12534
rect 4566 12470 4630 12534
rect 4647 12470 4711 12534
rect 4728 12470 4792 12534
rect 4809 12470 4873 12534
rect 105 12388 169 12452
rect 187 12388 251 12452
rect 269 12388 333 12452
rect 351 12388 415 12452
rect 433 12388 497 12452
rect 515 12388 579 12452
rect 597 12388 661 12452
rect 678 12388 742 12452
rect 759 12388 823 12452
rect 840 12388 904 12452
rect 921 12388 985 12452
rect 1002 12388 1066 12452
rect 1083 12388 1147 12452
rect 1164 12388 1228 12452
rect 1245 12388 1309 12452
rect 1326 12388 1390 12452
rect 1407 12388 1471 12452
rect 1488 12388 1552 12452
rect 1569 12388 1633 12452
rect 1650 12388 1714 12452
rect 1731 12388 1795 12452
rect 1812 12388 1876 12452
rect 1893 12388 1957 12452
rect 1974 12388 2038 12452
rect 2055 12388 2119 12452
rect 2136 12388 2200 12452
rect 2217 12388 2281 12452
rect 2298 12388 2362 12452
rect 2379 12388 2443 12452
rect 2460 12388 2524 12452
rect 2541 12388 2605 12452
rect 2622 12388 2686 12452
rect 2703 12388 2767 12452
rect 2784 12388 2848 12452
rect 2865 12388 2929 12452
rect 2946 12388 3010 12452
rect 3027 12388 3091 12452
rect 3108 12388 3172 12452
rect 3189 12388 3253 12452
rect 3270 12388 3334 12452
rect 3351 12388 3415 12452
rect 3432 12388 3496 12452
rect 3513 12388 3577 12452
rect 3594 12388 3658 12452
rect 3675 12388 3739 12452
rect 3756 12388 3820 12452
rect 3837 12388 3901 12452
rect 3918 12388 3982 12452
rect 3999 12388 4063 12452
rect 4080 12388 4144 12452
rect 4161 12388 4225 12452
rect 4242 12388 4306 12452
rect 4323 12388 4387 12452
rect 4404 12388 4468 12452
rect 4485 12388 4549 12452
rect 4566 12388 4630 12452
rect 4647 12388 4711 12452
rect 4728 12388 4792 12452
rect 4809 12388 4873 12452
rect 105 12306 169 12370
rect 187 12306 251 12370
rect 269 12306 333 12370
rect 351 12306 415 12370
rect 433 12306 497 12370
rect 515 12306 579 12370
rect 597 12306 661 12370
rect 678 12306 742 12370
rect 759 12306 823 12370
rect 840 12306 904 12370
rect 921 12306 985 12370
rect 1002 12306 1066 12370
rect 1083 12306 1147 12370
rect 1164 12306 1228 12370
rect 1245 12306 1309 12370
rect 1326 12306 1390 12370
rect 1407 12306 1471 12370
rect 1488 12306 1552 12370
rect 1569 12306 1633 12370
rect 1650 12306 1714 12370
rect 1731 12306 1795 12370
rect 1812 12306 1876 12370
rect 1893 12306 1957 12370
rect 1974 12306 2038 12370
rect 2055 12306 2119 12370
rect 2136 12306 2200 12370
rect 2217 12306 2281 12370
rect 2298 12306 2362 12370
rect 2379 12306 2443 12370
rect 2460 12306 2524 12370
rect 2541 12306 2605 12370
rect 2622 12306 2686 12370
rect 2703 12306 2767 12370
rect 2784 12306 2848 12370
rect 2865 12306 2929 12370
rect 2946 12306 3010 12370
rect 3027 12306 3091 12370
rect 3108 12306 3172 12370
rect 3189 12306 3253 12370
rect 3270 12306 3334 12370
rect 3351 12306 3415 12370
rect 3432 12306 3496 12370
rect 3513 12306 3577 12370
rect 3594 12306 3658 12370
rect 3675 12306 3739 12370
rect 3756 12306 3820 12370
rect 3837 12306 3901 12370
rect 3918 12306 3982 12370
rect 3999 12306 4063 12370
rect 4080 12306 4144 12370
rect 4161 12306 4225 12370
rect 4242 12306 4306 12370
rect 4323 12306 4387 12370
rect 4404 12306 4468 12370
rect 4485 12306 4549 12370
rect 4566 12306 4630 12370
rect 4647 12306 4711 12370
rect 4728 12306 4792 12370
rect 4809 12306 4873 12370
rect 105 12224 169 12288
rect 187 12224 251 12288
rect 269 12224 333 12288
rect 351 12224 415 12288
rect 433 12224 497 12288
rect 515 12224 579 12288
rect 597 12224 661 12288
rect 678 12224 742 12288
rect 759 12224 823 12288
rect 840 12224 904 12288
rect 921 12224 985 12288
rect 1002 12224 1066 12288
rect 1083 12224 1147 12288
rect 1164 12224 1228 12288
rect 1245 12224 1309 12288
rect 1326 12224 1390 12288
rect 1407 12224 1471 12288
rect 1488 12224 1552 12288
rect 1569 12224 1633 12288
rect 1650 12224 1714 12288
rect 1731 12224 1795 12288
rect 1812 12224 1876 12288
rect 1893 12224 1957 12288
rect 1974 12224 2038 12288
rect 2055 12224 2119 12288
rect 2136 12224 2200 12288
rect 2217 12224 2281 12288
rect 2298 12224 2362 12288
rect 2379 12224 2443 12288
rect 2460 12224 2524 12288
rect 2541 12224 2605 12288
rect 2622 12224 2686 12288
rect 2703 12224 2767 12288
rect 2784 12224 2848 12288
rect 2865 12224 2929 12288
rect 2946 12224 3010 12288
rect 3027 12224 3091 12288
rect 3108 12224 3172 12288
rect 3189 12224 3253 12288
rect 3270 12224 3334 12288
rect 3351 12224 3415 12288
rect 3432 12224 3496 12288
rect 3513 12224 3577 12288
rect 3594 12224 3658 12288
rect 3675 12224 3739 12288
rect 3756 12224 3820 12288
rect 3837 12224 3901 12288
rect 3918 12224 3982 12288
rect 3999 12224 4063 12288
rect 4080 12224 4144 12288
rect 4161 12224 4225 12288
rect 4242 12224 4306 12288
rect 4323 12224 4387 12288
rect 4404 12224 4468 12288
rect 4485 12224 4549 12288
rect 4566 12224 4630 12288
rect 4647 12224 4711 12288
rect 4728 12224 4792 12288
rect 4809 12224 4873 12288
rect 105 12142 169 12206
rect 187 12142 251 12206
rect 269 12142 333 12206
rect 351 12142 415 12206
rect 433 12142 497 12206
rect 515 12142 579 12206
rect 597 12142 661 12206
rect 678 12142 742 12206
rect 759 12142 823 12206
rect 840 12142 904 12206
rect 921 12142 985 12206
rect 1002 12142 1066 12206
rect 1083 12142 1147 12206
rect 1164 12142 1228 12206
rect 1245 12142 1309 12206
rect 1326 12142 1390 12206
rect 1407 12142 1471 12206
rect 1488 12142 1552 12206
rect 1569 12142 1633 12206
rect 1650 12142 1714 12206
rect 1731 12142 1795 12206
rect 1812 12142 1876 12206
rect 1893 12142 1957 12206
rect 1974 12142 2038 12206
rect 2055 12142 2119 12206
rect 2136 12142 2200 12206
rect 2217 12142 2281 12206
rect 2298 12142 2362 12206
rect 2379 12142 2443 12206
rect 2460 12142 2524 12206
rect 2541 12142 2605 12206
rect 2622 12142 2686 12206
rect 2703 12142 2767 12206
rect 2784 12142 2848 12206
rect 2865 12142 2929 12206
rect 2946 12142 3010 12206
rect 3027 12142 3091 12206
rect 3108 12142 3172 12206
rect 3189 12142 3253 12206
rect 3270 12142 3334 12206
rect 3351 12142 3415 12206
rect 3432 12142 3496 12206
rect 3513 12142 3577 12206
rect 3594 12142 3658 12206
rect 3675 12142 3739 12206
rect 3756 12142 3820 12206
rect 3837 12142 3901 12206
rect 3918 12142 3982 12206
rect 3999 12142 4063 12206
rect 4080 12142 4144 12206
rect 4161 12142 4225 12206
rect 4242 12142 4306 12206
rect 4323 12142 4387 12206
rect 4404 12142 4468 12206
rect 4485 12142 4549 12206
rect 4566 12142 4630 12206
rect 4647 12142 4711 12206
rect 4728 12142 4792 12206
rect 4809 12142 4873 12206
rect 105 12060 169 12124
rect 187 12060 251 12124
rect 269 12060 333 12124
rect 351 12060 415 12124
rect 433 12060 497 12124
rect 515 12060 579 12124
rect 597 12060 661 12124
rect 678 12060 742 12124
rect 759 12060 823 12124
rect 840 12060 904 12124
rect 921 12060 985 12124
rect 1002 12060 1066 12124
rect 1083 12060 1147 12124
rect 1164 12060 1228 12124
rect 1245 12060 1309 12124
rect 1326 12060 1390 12124
rect 1407 12060 1471 12124
rect 1488 12060 1552 12124
rect 1569 12060 1633 12124
rect 1650 12060 1714 12124
rect 1731 12060 1795 12124
rect 1812 12060 1876 12124
rect 1893 12060 1957 12124
rect 1974 12060 2038 12124
rect 2055 12060 2119 12124
rect 2136 12060 2200 12124
rect 2217 12060 2281 12124
rect 2298 12060 2362 12124
rect 2379 12060 2443 12124
rect 2460 12060 2524 12124
rect 2541 12060 2605 12124
rect 2622 12060 2686 12124
rect 2703 12060 2767 12124
rect 2784 12060 2848 12124
rect 2865 12060 2929 12124
rect 2946 12060 3010 12124
rect 3027 12060 3091 12124
rect 3108 12060 3172 12124
rect 3189 12060 3253 12124
rect 3270 12060 3334 12124
rect 3351 12060 3415 12124
rect 3432 12060 3496 12124
rect 3513 12060 3577 12124
rect 3594 12060 3658 12124
rect 3675 12060 3739 12124
rect 3756 12060 3820 12124
rect 3837 12060 3901 12124
rect 3918 12060 3982 12124
rect 3999 12060 4063 12124
rect 4080 12060 4144 12124
rect 4161 12060 4225 12124
rect 4242 12060 4306 12124
rect 4323 12060 4387 12124
rect 4404 12060 4468 12124
rect 4485 12060 4549 12124
rect 4566 12060 4630 12124
rect 4647 12060 4711 12124
rect 4728 12060 4792 12124
rect 4809 12060 4873 12124
rect 105 11978 169 12042
rect 187 11978 251 12042
rect 269 11978 333 12042
rect 351 11978 415 12042
rect 433 11978 497 12042
rect 515 11978 579 12042
rect 597 11978 661 12042
rect 678 11978 742 12042
rect 759 11978 823 12042
rect 840 11978 904 12042
rect 921 11978 985 12042
rect 1002 11978 1066 12042
rect 1083 11978 1147 12042
rect 1164 11978 1228 12042
rect 1245 11978 1309 12042
rect 1326 11978 1390 12042
rect 1407 11978 1471 12042
rect 1488 11978 1552 12042
rect 1569 11978 1633 12042
rect 1650 11978 1714 12042
rect 1731 11978 1795 12042
rect 1812 11978 1876 12042
rect 1893 11978 1957 12042
rect 1974 11978 2038 12042
rect 2055 11978 2119 12042
rect 2136 11978 2200 12042
rect 2217 11978 2281 12042
rect 2298 11978 2362 12042
rect 2379 11978 2443 12042
rect 2460 11978 2524 12042
rect 2541 11978 2605 12042
rect 2622 11978 2686 12042
rect 2703 11978 2767 12042
rect 2784 11978 2848 12042
rect 2865 11978 2929 12042
rect 2946 11978 3010 12042
rect 3027 11978 3091 12042
rect 3108 11978 3172 12042
rect 3189 11978 3253 12042
rect 3270 11978 3334 12042
rect 3351 11978 3415 12042
rect 3432 11978 3496 12042
rect 3513 11978 3577 12042
rect 3594 11978 3658 12042
rect 3675 11978 3739 12042
rect 3756 11978 3820 12042
rect 3837 11978 3901 12042
rect 3918 11978 3982 12042
rect 3999 11978 4063 12042
rect 4080 11978 4144 12042
rect 4161 11978 4225 12042
rect 4242 11978 4306 12042
rect 4323 11978 4387 12042
rect 4404 11978 4468 12042
rect 4485 11978 4549 12042
rect 4566 11978 4630 12042
rect 4647 11978 4711 12042
rect 4728 11978 4792 12042
rect 4809 11978 4873 12042
rect 105 11896 169 11960
rect 187 11896 251 11960
rect 269 11896 333 11960
rect 351 11896 415 11960
rect 433 11896 497 11960
rect 515 11896 579 11960
rect 597 11896 661 11960
rect 678 11896 742 11960
rect 759 11896 823 11960
rect 840 11896 904 11960
rect 921 11896 985 11960
rect 1002 11896 1066 11960
rect 1083 11896 1147 11960
rect 1164 11896 1228 11960
rect 1245 11896 1309 11960
rect 1326 11896 1390 11960
rect 1407 11896 1471 11960
rect 1488 11896 1552 11960
rect 1569 11896 1633 11960
rect 1650 11896 1714 11960
rect 1731 11896 1795 11960
rect 1812 11896 1876 11960
rect 1893 11896 1957 11960
rect 1974 11896 2038 11960
rect 2055 11896 2119 11960
rect 2136 11896 2200 11960
rect 2217 11896 2281 11960
rect 2298 11896 2362 11960
rect 2379 11896 2443 11960
rect 2460 11896 2524 11960
rect 2541 11896 2605 11960
rect 2622 11896 2686 11960
rect 2703 11896 2767 11960
rect 2784 11896 2848 11960
rect 2865 11896 2929 11960
rect 2946 11896 3010 11960
rect 3027 11896 3091 11960
rect 3108 11896 3172 11960
rect 3189 11896 3253 11960
rect 3270 11896 3334 11960
rect 3351 11896 3415 11960
rect 3432 11896 3496 11960
rect 3513 11896 3577 11960
rect 3594 11896 3658 11960
rect 3675 11896 3739 11960
rect 3756 11896 3820 11960
rect 3837 11896 3901 11960
rect 3918 11896 3982 11960
rect 3999 11896 4063 11960
rect 4080 11896 4144 11960
rect 4161 11896 4225 11960
rect 4242 11896 4306 11960
rect 4323 11896 4387 11960
rect 4404 11896 4468 11960
rect 4485 11896 4549 11960
rect 4566 11896 4630 11960
rect 4647 11896 4711 11960
rect 4728 11896 4792 11960
rect 4809 11896 4873 11960
rect 105 11814 169 11878
rect 187 11814 251 11878
rect 269 11814 333 11878
rect 351 11814 415 11878
rect 433 11814 497 11878
rect 515 11814 579 11878
rect 597 11814 661 11878
rect 678 11814 742 11878
rect 759 11814 823 11878
rect 840 11814 904 11878
rect 921 11814 985 11878
rect 1002 11814 1066 11878
rect 1083 11814 1147 11878
rect 1164 11814 1228 11878
rect 1245 11814 1309 11878
rect 1326 11814 1390 11878
rect 1407 11814 1471 11878
rect 1488 11814 1552 11878
rect 1569 11814 1633 11878
rect 1650 11814 1714 11878
rect 1731 11814 1795 11878
rect 1812 11814 1876 11878
rect 1893 11814 1957 11878
rect 1974 11814 2038 11878
rect 2055 11814 2119 11878
rect 2136 11814 2200 11878
rect 2217 11814 2281 11878
rect 2298 11814 2362 11878
rect 2379 11814 2443 11878
rect 2460 11814 2524 11878
rect 2541 11814 2605 11878
rect 2622 11814 2686 11878
rect 2703 11814 2767 11878
rect 2784 11814 2848 11878
rect 2865 11814 2929 11878
rect 2946 11814 3010 11878
rect 3027 11814 3091 11878
rect 3108 11814 3172 11878
rect 3189 11814 3253 11878
rect 3270 11814 3334 11878
rect 3351 11814 3415 11878
rect 3432 11814 3496 11878
rect 3513 11814 3577 11878
rect 3594 11814 3658 11878
rect 3675 11814 3739 11878
rect 3756 11814 3820 11878
rect 3837 11814 3901 11878
rect 3918 11814 3982 11878
rect 3999 11814 4063 11878
rect 4080 11814 4144 11878
rect 4161 11814 4225 11878
rect 4242 11814 4306 11878
rect 4323 11814 4387 11878
rect 4404 11814 4468 11878
rect 4485 11814 4549 11878
rect 4566 11814 4630 11878
rect 4647 11814 4711 11878
rect 4728 11814 4792 11878
rect 4809 11814 4873 11878
rect 105 11732 169 11796
rect 187 11732 251 11796
rect 269 11732 333 11796
rect 351 11732 415 11796
rect 433 11732 497 11796
rect 515 11732 579 11796
rect 597 11732 661 11796
rect 678 11732 742 11796
rect 759 11732 823 11796
rect 840 11732 904 11796
rect 921 11732 985 11796
rect 1002 11732 1066 11796
rect 1083 11732 1147 11796
rect 1164 11732 1228 11796
rect 1245 11732 1309 11796
rect 1326 11732 1390 11796
rect 1407 11732 1471 11796
rect 1488 11732 1552 11796
rect 1569 11732 1633 11796
rect 1650 11732 1714 11796
rect 1731 11732 1795 11796
rect 1812 11732 1876 11796
rect 1893 11732 1957 11796
rect 1974 11732 2038 11796
rect 2055 11732 2119 11796
rect 2136 11732 2200 11796
rect 2217 11732 2281 11796
rect 2298 11732 2362 11796
rect 2379 11732 2443 11796
rect 2460 11732 2524 11796
rect 2541 11732 2605 11796
rect 2622 11732 2686 11796
rect 2703 11732 2767 11796
rect 2784 11732 2848 11796
rect 2865 11732 2929 11796
rect 2946 11732 3010 11796
rect 3027 11732 3091 11796
rect 3108 11732 3172 11796
rect 3189 11732 3253 11796
rect 3270 11732 3334 11796
rect 3351 11732 3415 11796
rect 3432 11732 3496 11796
rect 3513 11732 3577 11796
rect 3594 11732 3658 11796
rect 3675 11732 3739 11796
rect 3756 11732 3820 11796
rect 3837 11732 3901 11796
rect 3918 11732 3982 11796
rect 3999 11732 4063 11796
rect 4080 11732 4144 11796
rect 4161 11732 4225 11796
rect 4242 11732 4306 11796
rect 4323 11732 4387 11796
rect 4404 11732 4468 11796
rect 4485 11732 4549 11796
rect 4566 11732 4630 11796
rect 4647 11732 4711 11796
rect 4728 11732 4792 11796
rect 4809 11732 4873 11796
rect 105 11650 169 11714
rect 187 11650 251 11714
rect 269 11650 333 11714
rect 351 11650 415 11714
rect 433 11650 497 11714
rect 515 11650 579 11714
rect 597 11650 661 11714
rect 678 11650 742 11714
rect 759 11650 823 11714
rect 840 11650 904 11714
rect 921 11650 985 11714
rect 1002 11650 1066 11714
rect 1083 11650 1147 11714
rect 1164 11650 1228 11714
rect 1245 11650 1309 11714
rect 1326 11650 1390 11714
rect 1407 11650 1471 11714
rect 1488 11650 1552 11714
rect 1569 11650 1633 11714
rect 1650 11650 1714 11714
rect 1731 11650 1795 11714
rect 1812 11650 1876 11714
rect 1893 11650 1957 11714
rect 1974 11650 2038 11714
rect 2055 11650 2119 11714
rect 2136 11650 2200 11714
rect 2217 11650 2281 11714
rect 2298 11650 2362 11714
rect 2379 11650 2443 11714
rect 2460 11650 2524 11714
rect 2541 11650 2605 11714
rect 2622 11650 2686 11714
rect 2703 11650 2767 11714
rect 2784 11650 2848 11714
rect 2865 11650 2929 11714
rect 2946 11650 3010 11714
rect 3027 11650 3091 11714
rect 3108 11650 3172 11714
rect 3189 11650 3253 11714
rect 3270 11650 3334 11714
rect 3351 11650 3415 11714
rect 3432 11650 3496 11714
rect 3513 11650 3577 11714
rect 3594 11650 3658 11714
rect 3675 11650 3739 11714
rect 3756 11650 3820 11714
rect 3837 11650 3901 11714
rect 3918 11650 3982 11714
rect 3999 11650 4063 11714
rect 4080 11650 4144 11714
rect 4161 11650 4225 11714
rect 4242 11650 4306 11714
rect 4323 11650 4387 11714
rect 4404 11650 4468 11714
rect 4485 11650 4549 11714
rect 4566 11650 4630 11714
rect 4647 11650 4711 11714
rect 4728 11650 4792 11714
rect 4809 11650 4873 11714
rect 10084 12470 10148 12534
rect 10166 12470 10230 12534
rect 10248 12470 10312 12534
rect 10330 12470 10394 12534
rect 10412 12470 10476 12534
rect 10494 12470 10558 12534
rect 10576 12470 10640 12534
rect 10657 12470 10721 12534
rect 10738 12470 10802 12534
rect 10819 12470 10883 12534
rect 10900 12470 10964 12534
rect 10981 12470 11045 12534
rect 11062 12470 11126 12534
rect 11143 12470 11207 12534
rect 11224 12470 11288 12534
rect 11305 12470 11369 12534
rect 11386 12470 11450 12534
rect 11467 12470 11531 12534
rect 11548 12470 11612 12534
rect 11629 12470 11693 12534
rect 11710 12470 11774 12534
rect 11791 12470 11855 12534
rect 11872 12470 11936 12534
rect 11953 12470 12017 12534
rect 12034 12470 12098 12534
rect 12115 12470 12179 12534
rect 12196 12470 12260 12534
rect 12277 12470 12341 12534
rect 12358 12470 12422 12534
rect 12439 12470 12503 12534
rect 12520 12470 12584 12534
rect 12601 12470 12665 12534
rect 12682 12470 12746 12534
rect 12763 12470 12827 12534
rect 12844 12470 12908 12534
rect 12925 12470 12989 12534
rect 13006 12470 13070 12534
rect 13087 12470 13151 12534
rect 13168 12470 13232 12534
rect 13249 12470 13313 12534
rect 13330 12470 13394 12534
rect 13411 12470 13475 12534
rect 13492 12470 13556 12534
rect 13573 12470 13637 12534
rect 13654 12470 13718 12534
rect 13735 12470 13799 12534
rect 13816 12470 13880 12534
rect 13897 12470 13961 12534
rect 13978 12470 14042 12534
rect 14059 12470 14123 12534
rect 14140 12470 14204 12534
rect 14221 12470 14285 12534
rect 14302 12470 14366 12534
rect 14383 12470 14447 12534
rect 14464 12470 14528 12534
rect 14545 12470 14609 12534
rect 14626 12470 14690 12534
rect 14707 12470 14771 12534
rect 14788 12470 14852 12534
rect 10084 12388 10148 12452
rect 10166 12388 10230 12452
rect 10248 12388 10312 12452
rect 10330 12388 10394 12452
rect 10412 12388 10476 12452
rect 10494 12388 10558 12452
rect 10576 12388 10640 12452
rect 10657 12388 10721 12452
rect 10738 12388 10802 12452
rect 10819 12388 10883 12452
rect 10900 12388 10964 12452
rect 10981 12388 11045 12452
rect 11062 12388 11126 12452
rect 11143 12388 11207 12452
rect 11224 12388 11288 12452
rect 11305 12388 11369 12452
rect 11386 12388 11450 12452
rect 11467 12388 11531 12452
rect 11548 12388 11612 12452
rect 11629 12388 11693 12452
rect 11710 12388 11774 12452
rect 11791 12388 11855 12452
rect 11872 12388 11936 12452
rect 11953 12388 12017 12452
rect 12034 12388 12098 12452
rect 12115 12388 12179 12452
rect 12196 12388 12260 12452
rect 12277 12388 12341 12452
rect 12358 12388 12422 12452
rect 12439 12388 12503 12452
rect 12520 12388 12584 12452
rect 12601 12388 12665 12452
rect 12682 12388 12746 12452
rect 12763 12388 12827 12452
rect 12844 12388 12908 12452
rect 12925 12388 12989 12452
rect 13006 12388 13070 12452
rect 13087 12388 13151 12452
rect 13168 12388 13232 12452
rect 13249 12388 13313 12452
rect 13330 12388 13394 12452
rect 13411 12388 13475 12452
rect 13492 12388 13556 12452
rect 13573 12388 13637 12452
rect 13654 12388 13718 12452
rect 13735 12388 13799 12452
rect 13816 12388 13880 12452
rect 13897 12388 13961 12452
rect 13978 12388 14042 12452
rect 14059 12388 14123 12452
rect 14140 12388 14204 12452
rect 14221 12388 14285 12452
rect 14302 12388 14366 12452
rect 14383 12388 14447 12452
rect 14464 12388 14528 12452
rect 14545 12388 14609 12452
rect 14626 12388 14690 12452
rect 14707 12388 14771 12452
rect 14788 12388 14852 12452
rect 10084 12306 10148 12370
rect 10166 12306 10230 12370
rect 10248 12306 10312 12370
rect 10330 12306 10394 12370
rect 10412 12306 10476 12370
rect 10494 12306 10558 12370
rect 10576 12306 10640 12370
rect 10657 12306 10721 12370
rect 10738 12306 10802 12370
rect 10819 12306 10883 12370
rect 10900 12306 10964 12370
rect 10981 12306 11045 12370
rect 11062 12306 11126 12370
rect 11143 12306 11207 12370
rect 11224 12306 11288 12370
rect 11305 12306 11369 12370
rect 11386 12306 11450 12370
rect 11467 12306 11531 12370
rect 11548 12306 11612 12370
rect 11629 12306 11693 12370
rect 11710 12306 11774 12370
rect 11791 12306 11855 12370
rect 11872 12306 11936 12370
rect 11953 12306 12017 12370
rect 12034 12306 12098 12370
rect 12115 12306 12179 12370
rect 12196 12306 12260 12370
rect 12277 12306 12341 12370
rect 12358 12306 12422 12370
rect 12439 12306 12503 12370
rect 12520 12306 12584 12370
rect 12601 12306 12665 12370
rect 12682 12306 12746 12370
rect 12763 12306 12827 12370
rect 12844 12306 12908 12370
rect 12925 12306 12989 12370
rect 13006 12306 13070 12370
rect 13087 12306 13151 12370
rect 13168 12306 13232 12370
rect 13249 12306 13313 12370
rect 13330 12306 13394 12370
rect 13411 12306 13475 12370
rect 13492 12306 13556 12370
rect 13573 12306 13637 12370
rect 13654 12306 13718 12370
rect 13735 12306 13799 12370
rect 13816 12306 13880 12370
rect 13897 12306 13961 12370
rect 13978 12306 14042 12370
rect 14059 12306 14123 12370
rect 14140 12306 14204 12370
rect 14221 12306 14285 12370
rect 14302 12306 14366 12370
rect 14383 12306 14447 12370
rect 14464 12306 14528 12370
rect 14545 12306 14609 12370
rect 14626 12306 14690 12370
rect 14707 12306 14771 12370
rect 14788 12306 14852 12370
rect 10084 12224 10148 12288
rect 10166 12224 10230 12288
rect 10248 12224 10312 12288
rect 10330 12224 10394 12288
rect 10412 12224 10476 12288
rect 10494 12224 10558 12288
rect 10576 12224 10640 12288
rect 10657 12224 10721 12288
rect 10738 12224 10802 12288
rect 10819 12224 10883 12288
rect 10900 12224 10964 12288
rect 10981 12224 11045 12288
rect 11062 12224 11126 12288
rect 11143 12224 11207 12288
rect 11224 12224 11288 12288
rect 11305 12224 11369 12288
rect 11386 12224 11450 12288
rect 11467 12224 11531 12288
rect 11548 12224 11612 12288
rect 11629 12224 11693 12288
rect 11710 12224 11774 12288
rect 11791 12224 11855 12288
rect 11872 12224 11936 12288
rect 11953 12224 12017 12288
rect 12034 12224 12098 12288
rect 12115 12224 12179 12288
rect 12196 12224 12260 12288
rect 12277 12224 12341 12288
rect 12358 12224 12422 12288
rect 12439 12224 12503 12288
rect 12520 12224 12584 12288
rect 12601 12224 12665 12288
rect 12682 12224 12746 12288
rect 12763 12224 12827 12288
rect 12844 12224 12908 12288
rect 12925 12224 12989 12288
rect 13006 12224 13070 12288
rect 13087 12224 13151 12288
rect 13168 12224 13232 12288
rect 13249 12224 13313 12288
rect 13330 12224 13394 12288
rect 13411 12224 13475 12288
rect 13492 12224 13556 12288
rect 13573 12224 13637 12288
rect 13654 12224 13718 12288
rect 13735 12224 13799 12288
rect 13816 12224 13880 12288
rect 13897 12224 13961 12288
rect 13978 12224 14042 12288
rect 14059 12224 14123 12288
rect 14140 12224 14204 12288
rect 14221 12224 14285 12288
rect 14302 12224 14366 12288
rect 14383 12224 14447 12288
rect 14464 12224 14528 12288
rect 14545 12224 14609 12288
rect 14626 12224 14690 12288
rect 14707 12224 14771 12288
rect 14788 12224 14852 12288
rect 10084 12142 10148 12206
rect 10166 12142 10230 12206
rect 10248 12142 10312 12206
rect 10330 12142 10394 12206
rect 10412 12142 10476 12206
rect 10494 12142 10558 12206
rect 10576 12142 10640 12206
rect 10657 12142 10721 12206
rect 10738 12142 10802 12206
rect 10819 12142 10883 12206
rect 10900 12142 10964 12206
rect 10981 12142 11045 12206
rect 11062 12142 11126 12206
rect 11143 12142 11207 12206
rect 11224 12142 11288 12206
rect 11305 12142 11369 12206
rect 11386 12142 11450 12206
rect 11467 12142 11531 12206
rect 11548 12142 11612 12206
rect 11629 12142 11693 12206
rect 11710 12142 11774 12206
rect 11791 12142 11855 12206
rect 11872 12142 11936 12206
rect 11953 12142 12017 12206
rect 12034 12142 12098 12206
rect 12115 12142 12179 12206
rect 12196 12142 12260 12206
rect 12277 12142 12341 12206
rect 12358 12142 12422 12206
rect 12439 12142 12503 12206
rect 12520 12142 12584 12206
rect 12601 12142 12665 12206
rect 12682 12142 12746 12206
rect 12763 12142 12827 12206
rect 12844 12142 12908 12206
rect 12925 12142 12989 12206
rect 13006 12142 13070 12206
rect 13087 12142 13151 12206
rect 13168 12142 13232 12206
rect 13249 12142 13313 12206
rect 13330 12142 13394 12206
rect 13411 12142 13475 12206
rect 13492 12142 13556 12206
rect 13573 12142 13637 12206
rect 13654 12142 13718 12206
rect 13735 12142 13799 12206
rect 13816 12142 13880 12206
rect 13897 12142 13961 12206
rect 13978 12142 14042 12206
rect 14059 12142 14123 12206
rect 14140 12142 14204 12206
rect 14221 12142 14285 12206
rect 14302 12142 14366 12206
rect 14383 12142 14447 12206
rect 14464 12142 14528 12206
rect 14545 12142 14609 12206
rect 14626 12142 14690 12206
rect 14707 12142 14771 12206
rect 14788 12142 14852 12206
rect 10084 12060 10148 12124
rect 10166 12060 10230 12124
rect 10248 12060 10312 12124
rect 10330 12060 10394 12124
rect 10412 12060 10476 12124
rect 10494 12060 10558 12124
rect 10576 12060 10640 12124
rect 10657 12060 10721 12124
rect 10738 12060 10802 12124
rect 10819 12060 10883 12124
rect 10900 12060 10964 12124
rect 10981 12060 11045 12124
rect 11062 12060 11126 12124
rect 11143 12060 11207 12124
rect 11224 12060 11288 12124
rect 11305 12060 11369 12124
rect 11386 12060 11450 12124
rect 11467 12060 11531 12124
rect 11548 12060 11612 12124
rect 11629 12060 11693 12124
rect 11710 12060 11774 12124
rect 11791 12060 11855 12124
rect 11872 12060 11936 12124
rect 11953 12060 12017 12124
rect 12034 12060 12098 12124
rect 12115 12060 12179 12124
rect 12196 12060 12260 12124
rect 12277 12060 12341 12124
rect 12358 12060 12422 12124
rect 12439 12060 12503 12124
rect 12520 12060 12584 12124
rect 12601 12060 12665 12124
rect 12682 12060 12746 12124
rect 12763 12060 12827 12124
rect 12844 12060 12908 12124
rect 12925 12060 12989 12124
rect 13006 12060 13070 12124
rect 13087 12060 13151 12124
rect 13168 12060 13232 12124
rect 13249 12060 13313 12124
rect 13330 12060 13394 12124
rect 13411 12060 13475 12124
rect 13492 12060 13556 12124
rect 13573 12060 13637 12124
rect 13654 12060 13718 12124
rect 13735 12060 13799 12124
rect 13816 12060 13880 12124
rect 13897 12060 13961 12124
rect 13978 12060 14042 12124
rect 14059 12060 14123 12124
rect 14140 12060 14204 12124
rect 14221 12060 14285 12124
rect 14302 12060 14366 12124
rect 14383 12060 14447 12124
rect 14464 12060 14528 12124
rect 14545 12060 14609 12124
rect 14626 12060 14690 12124
rect 14707 12060 14771 12124
rect 14788 12060 14852 12124
rect 10084 11978 10148 12042
rect 10166 11978 10230 12042
rect 10248 11978 10312 12042
rect 10330 11978 10394 12042
rect 10412 11978 10476 12042
rect 10494 11978 10558 12042
rect 10576 11978 10640 12042
rect 10657 11978 10721 12042
rect 10738 11978 10802 12042
rect 10819 11978 10883 12042
rect 10900 11978 10964 12042
rect 10981 11978 11045 12042
rect 11062 11978 11126 12042
rect 11143 11978 11207 12042
rect 11224 11978 11288 12042
rect 11305 11978 11369 12042
rect 11386 11978 11450 12042
rect 11467 11978 11531 12042
rect 11548 11978 11612 12042
rect 11629 11978 11693 12042
rect 11710 11978 11774 12042
rect 11791 11978 11855 12042
rect 11872 11978 11936 12042
rect 11953 11978 12017 12042
rect 12034 11978 12098 12042
rect 12115 11978 12179 12042
rect 12196 11978 12260 12042
rect 12277 11978 12341 12042
rect 12358 11978 12422 12042
rect 12439 11978 12503 12042
rect 12520 11978 12584 12042
rect 12601 11978 12665 12042
rect 12682 11978 12746 12042
rect 12763 11978 12827 12042
rect 12844 11978 12908 12042
rect 12925 11978 12989 12042
rect 13006 11978 13070 12042
rect 13087 11978 13151 12042
rect 13168 11978 13232 12042
rect 13249 11978 13313 12042
rect 13330 11978 13394 12042
rect 13411 11978 13475 12042
rect 13492 11978 13556 12042
rect 13573 11978 13637 12042
rect 13654 11978 13718 12042
rect 13735 11978 13799 12042
rect 13816 11978 13880 12042
rect 13897 11978 13961 12042
rect 13978 11978 14042 12042
rect 14059 11978 14123 12042
rect 14140 11978 14204 12042
rect 14221 11978 14285 12042
rect 14302 11978 14366 12042
rect 14383 11978 14447 12042
rect 14464 11978 14528 12042
rect 14545 11978 14609 12042
rect 14626 11978 14690 12042
rect 14707 11978 14771 12042
rect 14788 11978 14852 12042
rect 10084 11896 10148 11960
rect 10166 11896 10230 11960
rect 10248 11896 10312 11960
rect 10330 11896 10394 11960
rect 10412 11896 10476 11960
rect 10494 11896 10558 11960
rect 10576 11896 10640 11960
rect 10657 11896 10721 11960
rect 10738 11896 10802 11960
rect 10819 11896 10883 11960
rect 10900 11896 10964 11960
rect 10981 11896 11045 11960
rect 11062 11896 11126 11960
rect 11143 11896 11207 11960
rect 11224 11896 11288 11960
rect 11305 11896 11369 11960
rect 11386 11896 11450 11960
rect 11467 11896 11531 11960
rect 11548 11896 11612 11960
rect 11629 11896 11693 11960
rect 11710 11896 11774 11960
rect 11791 11896 11855 11960
rect 11872 11896 11936 11960
rect 11953 11896 12017 11960
rect 12034 11896 12098 11960
rect 12115 11896 12179 11960
rect 12196 11896 12260 11960
rect 12277 11896 12341 11960
rect 12358 11896 12422 11960
rect 12439 11896 12503 11960
rect 12520 11896 12584 11960
rect 12601 11896 12665 11960
rect 12682 11896 12746 11960
rect 12763 11896 12827 11960
rect 12844 11896 12908 11960
rect 12925 11896 12989 11960
rect 13006 11896 13070 11960
rect 13087 11896 13151 11960
rect 13168 11896 13232 11960
rect 13249 11896 13313 11960
rect 13330 11896 13394 11960
rect 13411 11896 13475 11960
rect 13492 11896 13556 11960
rect 13573 11896 13637 11960
rect 13654 11896 13718 11960
rect 13735 11896 13799 11960
rect 13816 11896 13880 11960
rect 13897 11896 13961 11960
rect 13978 11896 14042 11960
rect 14059 11896 14123 11960
rect 14140 11896 14204 11960
rect 14221 11896 14285 11960
rect 14302 11896 14366 11960
rect 14383 11896 14447 11960
rect 14464 11896 14528 11960
rect 14545 11896 14609 11960
rect 14626 11896 14690 11960
rect 14707 11896 14771 11960
rect 14788 11896 14852 11960
rect 10084 11814 10148 11878
rect 10166 11814 10230 11878
rect 10248 11814 10312 11878
rect 10330 11814 10394 11878
rect 10412 11814 10476 11878
rect 10494 11814 10558 11878
rect 10576 11814 10640 11878
rect 10657 11814 10721 11878
rect 10738 11814 10802 11878
rect 10819 11814 10883 11878
rect 10900 11814 10964 11878
rect 10981 11814 11045 11878
rect 11062 11814 11126 11878
rect 11143 11814 11207 11878
rect 11224 11814 11288 11878
rect 11305 11814 11369 11878
rect 11386 11814 11450 11878
rect 11467 11814 11531 11878
rect 11548 11814 11612 11878
rect 11629 11814 11693 11878
rect 11710 11814 11774 11878
rect 11791 11814 11855 11878
rect 11872 11814 11936 11878
rect 11953 11814 12017 11878
rect 12034 11814 12098 11878
rect 12115 11814 12179 11878
rect 12196 11814 12260 11878
rect 12277 11814 12341 11878
rect 12358 11814 12422 11878
rect 12439 11814 12503 11878
rect 12520 11814 12584 11878
rect 12601 11814 12665 11878
rect 12682 11814 12746 11878
rect 12763 11814 12827 11878
rect 12844 11814 12908 11878
rect 12925 11814 12989 11878
rect 13006 11814 13070 11878
rect 13087 11814 13151 11878
rect 13168 11814 13232 11878
rect 13249 11814 13313 11878
rect 13330 11814 13394 11878
rect 13411 11814 13475 11878
rect 13492 11814 13556 11878
rect 13573 11814 13637 11878
rect 13654 11814 13718 11878
rect 13735 11814 13799 11878
rect 13816 11814 13880 11878
rect 13897 11814 13961 11878
rect 13978 11814 14042 11878
rect 14059 11814 14123 11878
rect 14140 11814 14204 11878
rect 14221 11814 14285 11878
rect 14302 11814 14366 11878
rect 14383 11814 14447 11878
rect 14464 11814 14528 11878
rect 14545 11814 14609 11878
rect 14626 11814 14690 11878
rect 14707 11814 14771 11878
rect 14788 11814 14852 11878
rect 10084 11732 10148 11796
rect 10166 11732 10230 11796
rect 10248 11732 10312 11796
rect 10330 11732 10394 11796
rect 10412 11732 10476 11796
rect 10494 11732 10558 11796
rect 10576 11732 10640 11796
rect 10657 11732 10721 11796
rect 10738 11732 10802 11796
rect 10819 11732 10883 11796
rect 10900 11732 10964 11796
rect 10981 11732 11045 11796
rect 11062 11732 11126 11796
rect 11143 11732 11207 11796
rect 11224 11732 11288 11796
rect 11305 11732 11369 11796
rect 11386 11732 11450 11796
rect 11467 11732 11531 11796
rect 11548 11732 11612 11796
rect 11629 11732 11693 11796
rect 11710 11732 11774 11796
rect 11791 11732 11855 11796
rect 11872 11732 11936 11796
rect 11953 11732 12017 11796
rect 12034 11732 12098 11796
rect 12115 11732 12179 11796
rect 12196 11732 12260 11796
rect 12277 11732 12341 11796
rect 12358 11732 12422 11796
rect 12439 11732 12503 11796
rect 12520 11732 12584 11796
rect 12601 11732 12665 11796
rect 12682 11732 12746 11796
rect 12763 11732 12827 11796
rect 12844 11732 12908 11796
rect 12925 11732 12989 11796
rect 13006 11732 13070 11796
rect 13087 11732 13151 11796
rect 13168 11732 13232 11796
rect 13249 11732 13313 11796
rect 13330 11732 13394 11796
rect 13411 11732 13475 11796
rect 13492 11732 13556 11796
rect 13573 11732 13637 11796
rect 13654 11732 13718 11796
rect 13735 11732 13799 11796
rect 13816 11732 13880 11796
rect 13897 11732 13961 11796
rect 13978 11732 14042 11796
rect 14059 11732 14123 11796
rect 14140 11732 14204 11796
rect 14221 11732 14285 11796
rect 14302 11732 14366 11796
rect 14383 11732 14447 11796
rect 14464 11732 14528 11796
rect 14545 11732 14609 11796
rect 14626 11732 14690 11796
rect 14707 11732 14771 11796
rect 14788 11732 14852 11796
rect 10084 11650 10148 11714
rect 10166 11650 10230 11714
rect 10248 11650 10312 11714
rect 10330 11650 10394 11714
rect 10412 11650 10476 11714
rect 10494 11650 10558 11714
rect 10576 11650 10640 11714
rect 10657 11650 10721 11714
rect 10738 11650 10802 11714
rect 10819 11650 10883 11714
rect 10900 11650 10964 11714
rect 10981 11650 11045 11714
rect 11062 11650 11126 11714
rect 11143 11650 11207 11714
rect 11224 11650 11288 11714
rect 11305 11650 11369 11714
rect 11386 11650 11450 11714
rect 11467 11650 11531 11714
rect 11548 11650 11612 11714
rect 11629 11650 11693 11714
rect 11710 11650 11774 11714
rect 11791 11650 11855 11714
rect 11872 11650 11936 11714
rect 11953 11650 12017 11714
rect 12034 11650 12098 11714
rect 12115 11650 12179 11714
rect 12196 11650 12260 11714
rect 12277 11650 12341 11714
rect 12358 11650 12422 11714
rect 12439 11650 12503 11714
rect 12520 11650 12584 11714
rect 12601 11650 12665 11714
rect 12682 11650 12746 11714
rect 12763 11650 12827 11714
rect 12844 11650 12908 11714
rect 12925 11650 12989 11714
rect 13006 11650 13070 11714
rect 13087 11650 13151 11714
rect 13168 11650 13232 11714
rect 13249 11650 13313 11714
rect 13330 11650 13394 11714
rect 13411 11650 13475 11714
rect 13492 11650 13556 11714
rect 13573 11650 13637 11714
rect 13654 11650 13718 11714
rect 13735 11650 13799 11714
rect 13816 11650 13880 11714
rect 13897 11650 13961 11714
rect 13978 11650 14042 11714
rect 14059 11650 14123 11714
rect 14140 11650 14204 11714
rect 14221 11650 14285 11714
rect 14302 11650 14366 11714
rect 14383 11650 14447 11714
rect 14464 11650 14528 11714
rect 14545 11650 14609 11714
rect 14626 11650 14690 11714
rect 14707 11650 14771 11714
rect 14788 11650 14852 11714
rect 105 6030 169 6094
rect 187 6030 251 6094
rect 269 6030 333 6094
rect 351 6030 415 6094
rect 433 6030 497 6094
rect 515 6030 579 6094
rect 597 6030 661 6094
rect 678 6030 742 6094
rect 759 6030 823 6094
rect 840 6030 904 6094
rect 921 6030 985 6094
rect 1002 6030 1066 6094
rect 1083 6030 1147 6094
rect 1164 6030 1228 6094
rect 1245 6030 1309 6094
rect 1326 6030 1390 6094
rect 1407 6030 1471 6094
rect 1488 6030 1552 6094
rect 1569 6030 1633 6094
rect 1650 6030 1714 6094
rect 1731 6030 1795 6094
rect 1812 6030 1876 6094
rect 1893 6030 1957 6094
rect 1974 6030 2038 6094
rect 2055 6030 2119 6094
rect 2136 6030 2200 6094
rect 2217 6030 2281 6094
rect 2298 6030 2362 6094
rect 2379 6030 2443 6094
rect 2460 6030 2524 6094
rect 2541 6030 2605 6094
rect 2622 6030 2686 6094
rect 2703 6030 2767 6094
rect 2784 6030 2848 6094
rect 2865 6030 2929 6094
rect 2946 6030 3010 6094
rect 3027 6030 3091 6094
rect 3108 6030 3172 6094
rect 3189 6030 3253 6094
rect 3270 6030 3334 6094
rect 3351 6030 3415 6094
rect 3432 6030 3496 6094
rect 3513 6030 3577 6094
rect 3594 6030 3658 6094
rect 3675 6030 3739 6094
rect 3756 6030 3820 6094
rect 3837 6030 3901 6094
rect 3918 6030 3982 6094
rect 3999 6030 4063 6094
rect 4080 6030 4144 6094
rect 4161 6030 4225 6094
rect 4242 6030 4306 6094
rect 4323 6030 4387 6094
rect 4404 6030 4468 6094
rect 4485 6030 4549 6094
rect 4566 6030 4630 6094
rect 4647 6030 4711 6094
rect 4728 6030 4792 6094
rect 4809 6030 4873 6094
rect 105 5944 169 6008
rect 187 5944 251 6008
rect 269 5944 333 6008
rect 351 5944 415 6008
rect 433 5944 497 6008
rect 515 5944 579 6008
rect 597 5944 661 6008
rect 678 5944 742 6008
rect 759 5944 823 6008
rect 840 5944 904 6008
rect 921 5944 985 6008
rect 1002 5944 1066 6008
rect 1083 5944 1147 6008
rect 1164 5944 1228 6008
rect 1245 5944 1309 6008
rect 1326 5944 1390 6008
rect 1407 5944 1471 6008
rect 1488 5944 1552 6008
rect 1569 5944 1633 6008
rect 1650 5944 1714 6008
rect 1731 5944 1795 6008
rect 1812 5944 1876 6008
rect 1893 5944 1957 6008
rect 1974 5944 2038 6008
rect 2055 5944 2119 6008
rect 2136 5944 2200 6008
rect 2217 5944 2281 6008
rect 2298 5944 2362 6008
rect 2379 5944 2443 6008
rect 2460 5944 2524 6008
rect 2541 5944 2605 6008
rect 2622 5944 2686 6008
rect 2703 5944 2767 6008
rect 2784 5944 2848 6008
rect 2865 5944 2929 6008
rect 2946 5944 3010 6008
rect 3027 5944 3091 6008
rect 3108 5944 3172 6008
rect 3189 5944 3253 6008
rect 3270 5944 3334 6008
rect 3351 5944 3415 6008
rect 3432 5944 3496 6008
rect 3513 5944 3577 6008
rect 3594 5944 3658 6008
rect 3675 5944 3739 6008
rect 3756 5944 3820 6008
rect 3837 5944 3901 6008
rect 3918 5944 3982 6008
rect 3999 5944 4063 6008
rect 4080 5944 4144 6008
rect 4161 5944 4225 6008
rect 4242 5944 4306 6008
rect 4323 5944 4387 6008
rect 4404 5944 4468 6008
rect 4485 5944 4549 6008
rect 4566 5944 4630 6008
rect 4647 5944 4711 6008
rect 4728 5944 4792 6008
rect 4809 5944 4873 6008
rect 105 5858 169 5922
rect 187 5858 251 5922
rect 269 5858 333 5922
rect 351 5858 415 5922
rect 433 5858 497 5922
rect 515 5858 579 5922
rect 597 5858 661 5922
rect 678 5858 742 5922
rect 759 5858 823 5922
rect 840 5858 904 5922
rect 921 5858 985 5922
rect 1002 5858 1066 5922
rect 1083 5858 1147 5922
rect 1164 5858 1228 5922
rect 1245 5858 1309 5922
rect 1326 5858 1390 5922
rect 1407 5858 1471 5922
rect 1488 5858 1552 5922
rect 1569 5858 1633 5922
rect 1650 5858 1714 5922
rect 1731 5858 1795 5922
rect 1812 5858 1876 5922
rect 1893 5858 1957 5922
rect 1974 5858 2038 5922
rect 2055 5858 2119 5922
rect 2136 5858 2200 5922
rect 2217 5858 2281 5922
rect 2298 5858 2362 5922
rect 2379 5858 2443 5922
rect 2460 5858 2524 5922
rect 2541 5858 2605 5922
rect 2622 5858 2686 5922
rect 2703 5858 2767 5922
rect 2784 5858 2848 5922
rect 2865 5858 2929 5922
rect 2946 5858 3010 5922
rect 3027 5858 3091 5922
rect 3108 5858 3172 5922
rect 3189 5858 3253 5922
rect 3270 5858 3334 5922
rect 3351 5858 3415 5922
rect 3432 5858 3496 5922
rect 3513 5858 3577 5922
rect 3594 5858 3658 5922
rect 3675 5858 3739 5922
rect 3756 5858 3820 5922
rect 3837 5858 3901 5922
rect 3918 5858 3982 5922
rect 3999 5858 4063 5922
rect 4080 5858 4144 5922
rect 4161 5858 4225 5922
rect 4242 5858 4306 5922
rect 4323 5858 4387 5922
rect 4404 5858 4468 5922
rect 4485 5858 4549 5922
rect 4566 5858 4630 5922
rect 4647 5858 4711 5922
rect 4728 5858 4792 5922
rect 4809 5858 4873 5922
rect 105 5772 169 5836
rect 187 5772 251 5836
rect 269 5772 333 5836
rect 351 5772 415 5836
rect 433 5772 497 5836
rect 515 5772 579 5836
rect 597 5772 661 5836
rect 678 5772 742 5836
rect 759 5772 823 5836
rect 840 5772 904 5836
rect 921 5772 985 5836
rect 1002 5772 1066 5836
rect 1083 5772 1147 5836
rect 1164 5772 1228 5836
rect 1245 5772 1309 5836
rect 1326 5772 1390 5836
rect 1407 5772 1471 5836
rect 1488 5772 1552 5836
rect 1569 5772 1633 5836
rect 1650 5772 1714 5836
rect 1731 5772 1795 5836
rect 1812 5772 1876 5836
rect 1893 5772 1957 5836
rect 1974 5772 2038 5836
rect 2055 5772 2119 5836
rect 2136 5772 2200 5836
rect 2217 5772 2281 5836
rect 2298 5772 2362 5836
rect 2379 5772 2443 5836
rect 2460 5772 2524 5836
rect 2541 5772 2605 5836
rect 2622 5772 2686 5836
rect 2703 5772 2767 5836
rect 2784 5772 2848 5836
rect 2865 5772 2929 5836
rect 2946 5772 3010 5836
rect 3027 5772 3091 5836
rect 3108 5772 3172 5836
rect 3189 5772 3253 5836
rect 3270 5772 3334 5836
rect 3351 5772 3415 5836
rect 3432 5772 3496 5836
rect 3513 5772 3577 5836
rect 3594 5772 3658 5836
rect 3675 5772 3739 5836
rect 3756 5772 3820 5836
rect 3837 5772 3901 5836
rect 3918 5772 3982 5836
rect 3999 5772 4063 5836
rect 4080 5772 4144 5836
rect 4161 5772 4225 5836
rect 4242 5772 4306 5836
rect 4323 5772 4387 5836
rect 4404 5772 4468 5836
rect 4485 5772 4549 5836
rect 4566 5772 4630 5836
rect 4647 5772 4711 5836
rect 4728 5772 4792 5836
rect 4809 5772 4873 5836
rect 105 5686 169 5750
rect 187 5686 251 5750
rect 269 5686 333 5750
rect 351 5686 415 5750
rect 433 5686 497 5750
rect 515 5686 579 5750
rect 597 5686 661 5750
rect 678 5686 742 5750
rect 759 5686 823 5750
rect 840 5686 904 5750
rect 921 5686 985 5750
rect 1002 5686 1066 5750
rect 1083 5686 1147 5750
rect 1164 5686 1228 5750
rect 1245 5686 1309 5750
rect 1326 5686 1390 5750
rect 1407 5686 1471 5750
rect 1488 5686 1552 5750
rect 1569 5686 1633 5750
rect 1650 5686 1714 5750
rect 1731 5686 1795 5750
rect 1812 5686 1876 5750
rect 1893 5686 1957 5750
rect 1974 5686 2038 5750
rect 2055 5686 2119 5750
rect 2136 5686 2200 5750
rect 2217 5686 2281 5750
rect 2298 5686 2362 5750
rect 2379 5686 2443 5750
rect 2460 5686 2524 5750
rect 2541 5686 2605 5750
rect 2622 5686 2686 5750
rect 2703 5686 2767 5750
rect 2784 5686 2848 5750
rect 2865 5686 2929 5750
rect 2946 5686 3010 5750
rect 3027 5686 3091 5750
rect 3108 5686 3172 5750
rect 3189 5686 3253 5750
rect 3270 5686 3334 5750
rect 3351 5686 3415 5750
rect 3432 5686 3496 5750
rect 3513 5686 3577 5750
rect 3594 5686 3658 5750
rect 3675 5686 3739 5750
rect 3756 5686 3820 5750
rect 3837 5686 3901 5750
rect 3918 5686 3982 5750
rect 3999 5686 4063 5750
rect 4080 5686 4144 5750
rect 4161 5686 4225 5750
rect 4242 5686 4306 5750
rect 4323 5686 4387 5750
rect 4404 5686 4468 5750
rect 4485 5686 4549 5750
rect 4566 5686 4630 5750
rect 4647 5686 4711 5750
rect 4728 5686 4792 5750
rect 4809 5686 4873 5750
rect 105 5600 169 5664
rect 187 5600 251 5664
rect 269 5600 333 5664
rect 351 5600 415 5664
rect 433 5600 497 5664
rect 515 5600 579 5664
rect 597 5600 661 5664
rect 678 5600 742 5664
rect 759 5600 823 5664
rect 840 5600 904 5664
rect 921 5600 985 5664
rect 1002 5600 1066 5664
rect 1083 5600 1147 5664
rect 1164 5600 1228 5664
rect 1245 5600 1309 5664
rect 1326 5600 1390 5664
rect 1407 5600 1471 5664
rect 1488 5600 1552 5664
rect 1569 5600 1633 5664
rect 1650 5600 1714 5664
rect 1731 5600 1795 5664
rect 1812 5600 1876 5664
rect 1893 5600 1957 5664
rect 1974 5600 2038 5664
rect 2055 5600 2119 5664
rect 2136 5600 2200 5664
rect 2217 5600 2281 5664
rect 2298 5600 2362 5664
rect 2379 5600 2443 5664
rect 2460 5600 2524 5664
rect 2541 5600 2605 5664
rect 2622 5600 2686 5664
rect 2703 5600 2767 5664
rect 2784 5600 2848 5664
rect 2865 5600 2929 5664
rect 2946 5600 3010 5664
rect 3027 5600 3091 5664
rect 3108 5600 3172 5664
rect 3189 5600 3253 5664
rect 3270 5600 3334 5664
rect 3351 5600 3415 5664
rect 3432 5600 3496 5664
rect 3513 5600 3577 5664
rect 3594 5600 3658 5664
rect 3675 5600 3739 5664
rect 3756 5600 3820 5664
rect 3837 5600 3901 5664
rect 3918 5600 3982 5664
rect 3999 5600 4063 5664
rect 4080 5600 4144 5664
rect 4161 5600 4225 5664
rect 4242 5600 4306 5664
rect 4323 5600 4387 5664
rect 4404 5600 4468 5664
rect 4485 5600 4549 5664
rect 4566 5600 4630 5664
rect 4647 5600 4711 5664
rect 4728 5600 4792 5664
rect 4809 5600 4873 5664
rect 105 5514 169 5578
rect 187 5514 251 5578
rect 269 5514 333 5578
rect 351 5514 415 5578
rect 433 5514 497 5578
rect 515 5514 579 5578
rect 597 5514 661 5578
rect 678 5514 742 5578
rect 759 5514 823 5578
rect 840 5514 904 5578
rect 921 5514 985 5578
rect 1002 5514 1066 5578
rect 1083 5514 1147 5578
rect 1164 5514 1228 5578
rect 1245 5514 1309 5578
rect 1326 5514 1390 5578
rect 1407 5514 1471 5578
rect 1488 5514 1552 5578
rect 1569 5514 1633 5578
rect 1650 5514 1714 5578
rect 1731 5514 1795 5578
rect 1812 5514 1876 5578
rect 1893 5514 1957 5578
rect 1974 5514 2038 5578
rect 2055 5514 2119 5578
rect 2136 5514 2200 5578
rect 2217 5514 2281 5578
rect 2298 5514 2362 5578
rect 2379 5514 2443 5578
rect 2460 5514 2524 5578
rect 2541 5514 2605 5578
rect 2622 5514 2686 5578
rect 2703 5514 2767 5578
rect 2784 5514 2848 5578
rect 2865 5514 2929 5578
rect 2946 5514 3010 5578
rect 3027 5514 3091 5578
rect 3108 5514 3172 5578
rect 3189 5514 3253 5578
rect 3270 5514 3334 5578
rect 3351 5514 3415 5578
rect 3432 5514 3496 5578
rect 3513 5514 3577 5578
rect 3594 5514 3658 5578
rect 3675 5514 3739 5578
rect 3756 5514 3820 5578
rect 3837 5514 3901 5578
rect 3918 5514 3982 5578
rect 3999 5514 4063 5578
rect 4080 5514 4144 5578
rect 4161 5514 4225 5578
rect 4242 5514 4306 5578
rect 4323 5514 4387 5578
rect 4404 5514 4468 5578
rect 4485 5514 4549 5578
rect 4566 5514 4630 5578
rect 4647 5514 4711 5578
rect 4728 5514 4792 5578
rect 4809 5514 4873 5578
rect 105 5428 169 5492
rect 187 5428 251 5492
rect 269 5428 333 5492
rect 351 5428 415 5492
rect 433 5428 497 5492
rect 515 5428 579 5492
rect 597 5428 661 5492
rect 678 5428 742 5492
rect 759 5428 823 5492
rect 840 5428 904 5492
rect 921 5428 985 5492
rect 1002 5428 1066 5492
rect 1083 5428 1147 5492
rect 1164 5428 1228 5492
rect 1245 5428 1309 5492
rect 1326 5428 1390 5492
rect 1407 5428 1471 5492
rect 1488 5428 1552 5492
rect 1569 5428 1633 5492
rect 1650 5428 1714 5492
rect 1731 5428 1795 5492
rect 1812 5428 1876 5492
rect 1893 5428 1957 5492
rect 1974 5428 2038 5492
rect 2055 5428 2119 5492
rect 2136 5428 2200 5492
rect 2217 5428 2281 5492
rect 2298 5428 2362 5492
rect 2379 5428 2443 5492
rect 2460 5428 2524 5492
rect 2541 5428 2605 5492
rect 2622 5428 2686 5492
rect 2703 5428 2767 5492
rect 2784 5428 2848 5492
rect 2865 5428 2929 5492
rect 2946 5428 3010 5492
rect 3027 5428 3091 5492
rect 3108 5428 3172 5492
rect 3189 5428 3253 5492
rect 3270 5428 3334 5492
rect 3351 5428 3415 5492
rect 3432 5428 3496 5492
rect 3513 5428 3577 5492
rect 3594 5428 3658 5492
rect 3675 5428 3739 5492
rect 3756 5428 3820 5492
rect 3837 5428 3901 5492
rect 3918 5428 3982 5492
rect 3999 5428 4063 5492
rect 4080 5428 4144 5492
rect 4161 5428 4225 5492
rect 4242 5428 4306 5492
rect 4323 5428 4387 5492
rect 4404 5428 4468 5492
rect 4485 5428 4549 5492
rect 4566 5428 4630 5492
rect 4647 5428 4711 5492
rect 4728 5428 4792 5492
rect 4809 5428 4873 5492
rect 105 5342 169 5406
rect 187 5342 251 5406
rect 269 5342 333 5406
rect 351 5342 415 5406
rect 433 5342 497 5406
rect 515 5342 579 5406
rect 597 5342 661 5406
rect 678 5342 742 5406
rect 759 5342 823 5406
rect 840 5342 904 5406
rect 921 5342 985 5406
rect 1002 5342 1066 5406
rect 1083 5342 1147 5406
rect 1164 5342 1228 5406
rect 1245 5342 1309 5406
rect 1326 5342 1390 5406
rect 1407 5342 1471 5406
rect 1488 5342 1552 5406
rect 1569 5342 1633 5406
rect 1650 5342 1714 5406
rect 1731 5342 1795 5406
rect 1812 5342 1876 5406
rect 1893 5342 1957 5406
rect 1974 5342 2038 5406
rect 2055 5342 2119 5406
rect 2136 5342 2200 5406
rect 2217 5342 2281 5406
rect 2298 5342 2362 5406
rect 2379 5342 2443 5406
rect 2460 5342 2524 5406
rect 2541 5342 2605 5406
rect 2622 5342 2686 5406
rect 2703 5342 2767 5406
rect 2784 5342 2848 5406
rect 2865 5342 2929 5406
rect 2946 5342 3010 5406
rect 3027 5342 3091 5406
rect 3108 5342 3172 5406
rect 3189 5342 3253 5406
rect 3270 5342 3334 5406
rect 3351 5342 3415 5406
rect 3432 5342 3496 5406
rect 3513 5342 3577 5406
rect 3594 5342 3658 5406
rect 3675 5342 3739 5406
rect 3756 5342 3820 5406
rect 3837 5342 3901 5406
rect 3918 5342 3982 5406
rect 3999 5342 4063 5406
rect 4080 5342 4144 5406
rect 4161 5342 4225 5406
rect 4242 5342 4306 5406
rect 4323 5342 4387 5406
rect 4404 5342 4468 5406
rect 4485 5342 4549 5406
rect 4566 5342 4630 5406
rect 4647 5342 4711 5406
rect 4728 5342 4792 5406
rect 4809 5342 4873 5406
rect 105 5256 169 5320
rect 187 5256 251 5320
rect 269 5256 333 5320
rect 351 5256 415 5320
rect 433 5256 497 5320
rect 515 5256 579 5320
rect 597 5256 661 5320
rect 678 5256 742 5320
rect 759 5256 823 5320
rect 840 5256 904 5320
rect 921 5256 985 5320
rect 1002 5256 1066 5320
rect 1083 5256 1147 5320
rect 1164 5256 1228 5320
rect 1245 5256 1309 5320
rect 1326 5256 1390 5320
rect 1407 5256 1471 5320
rect 1488 5256 1552 5320
rect 1569 5256 1633 5320
rect 1650 5256 1714 5320
rect 1731 5256 1795 5320
rect 1812 5256 1876 5320
rect 1893 5256 1957 5320
rect 1974 5256 2038 5320
rect 2055 5256 2119 5320
rect 2136 5256 2200 5320
rect 2217 5256 2281 5320
rect 2298 5256 2362 5320
rect 2379 5256 2443 5320
rect 2460 5256 2524 5320
rect 2541 5256 2605 5320
rect 2622 5256 2686 5320
rect 2703 5256 2767 5320
rect 2784 5256 2848 5320
rect 2865 5256 2929 5320
rect 2946 5256 3010 5320
rect 3027 5256 3091 5320
rect 3108 5256 3172 5320
rect 3189 5256 3253 5320
rect 3270 5256 3334 5320
rect 3351 5256 3415 5320
rect 3432 5256 3496 5320
rect 3513 5256 3577 5320
rect 3594 5256 3658 5320
rect 3675 5256 3739 5320
rect 3756 5256 3820 5320
rect 3837 5256 3901 5320
rect 3918 5256 3982 5320
rect 3999 5256 4063 5320
rect 4080 5256 4144 5320
rect 4161 5256 4225 5320
rect 4242 5256 4306 5320
rect 4323 5256 4387 5320
rect 4404 5256 4468 5320
rect 4485 5256 4549 5320
rect 4566 5256 4630 5320
rect 4647 5256 4711 5320
rect 4728 5256 4792 5320
rect 4809 5256 4873 5320
rect 105 5170 169 5234
rect 187 5170 251 5234
rect 269 5170 333 5234
rect 351 5170 415 5234
rect 433 5170 497 5234
rect 515 5170 579 5234
rect 597 5170 661 5234
rect 678 5170 742 5234
rect 759 5170 823 5234
rect 840 5170 904 5234
rect 921 5170 985 5234
rect 1002 5170 1066 5234
rect 1083 5170 1147 5234
rect 1164 5170 1228 5234
rect 1245 5170 1309 5234
rect 1326 5170 1390 5234
rect 1407 5170 1471 5234
rect 1488 5170 1552 5234
rect 1569 5170 1633 5234
rect 1650 5170 1714 5234
rect 1731 5170 1795 5234
rect 1812 5170 1876 5234
rect 1893 5170 1957 5234
rect 1974 5170 2038 5234
rect 2055 5170 2119 5234
rect 2136 5170 2200 5234
rect 2217 5170 2281 5234
rect 2298 5170 2362 5234
rect 2379 5170 2443 5234
rect 2460 5170 2524 5234
rect 2541 5170 2605 5234
rect 2622 5170 2686 5234
rect 2703 5170 2767 5234
rect 2784 5170 2848 5234
rect 2865 5170 2929 5234
rect 2946 5170 3010 5234
rect 3027 5170 3091 5234
rect 3108 5170 3172 5234
rect 3189 5170 3253 5234
rect 3270 5170 3334 5234
rect 3351 5170 3415 5234
rect 3432 5170 3496 5234
rect 3513 5170 3577 5234
rect 3594 5170 3658 5234
rect 3675 5170 3739 5234
rect 3756 5170 3820 5234
rect 3837 5170 3901 5234
rect 3918 5170 3982 5234
rect 3999 5170 4063 5234
rect 4080 5170 4144 5234
rect 4161 5170 4225 5234
rect 4242 5170 4306 5234
rect 4323 5170 4387 5234
rect 4404 5170 4468 5234
rect 4485 5170 4549 5234
rect 4566 5170 4630 5234
rect 4647 5170 4711 5234
rect 4728 5170 4792 5234
rect 4809 5170 4873 5234
rect 10084 6030 10148 6094
rect 10166 6030 10230 6094
rect 10248 6030 10312 6094
rect 10330 6030 10394 6094
rect 10412 6030 10476 6094
rect 10494 6030 10558 6094
rect 10576 6030 10640 6094
rect 10657 6030 10721 6094
rect 10738 6030 10802 6094
rect 10819 6030 10883 6094
rect 10900 6030 10964 6094
rect 10981 6030 11045 6094
rect 11062 6030 11126 6094
rect 11143 6030 11207 6094
rect 11224 6030 11288 6094
rect 11305 6030 11369 6094
rect 11386 6030 11450 6094
rect 11467 6030 11531 6094
rect 11548 6030 11612 6094
rect 11629 6030 11693 6094
rect 11710 6030 11774 6094
rect 11791 6030 11855 6094
rect 11872 6030 11936 6094
rect 11953 6030 12017 6094
rect 12034 6030 12098 6094
rect 12115 6030 12179 6094
rect 12196 6030 12260 6094
rect 12277 6030 12341 6094
rect 12358 6030 12422 6094
rect 12439 6030 12503 6094
rect 12520 6030 12584 6094
rect 12601 6030 12665 6094
rect 12682 6030 12746 6094
rect 12763 6030 12827 6094
rect 12844 6030 12908 6094
rect 12925 6030 12989 6094
rect 13006 6030 13070 6094
rect 13087 6030 13151 6094
rect 13168 6030 13232 6094
rect 13249 6030 13313 6094
rect 13330 6030 13394 6094
rect 13411 6030 13475 6094
rect 13492 6030 13556 6094
rect 13573 6030 13637 6094
rect 13654 6030 13718 6094
rect 13735 6030 13799 6094
rect 13816 6030 13880 6094
rect 13897 6030 13961 6094
rect 13978 6030 14042 6094
rect 14059 6030 14123 6094
rect 14140 6030 14204 6094
rect 14221 6030 14285 6094
rect 14302 6030 14366 6094
rect 14383 6030 14447 6094
rect 14464 6030 14528 6094
rect 14545 6030 14609 6094
rect 14626 6030 14690 6094
rect 14707 6030 14771 6094
rect 14788 6030 14852 6094
rect 10084 5944 10148 6008
rect 10166 5944 10230 6008
rect 10248 5944 10312 6008
rect 10330 5944 10394 6008
rect 10412 5944 10476 6008
rect 10494 5944 10558 6008
rect 10576 5944 10640 6008
rect 10657 5944 10721 6008
rect 10738 5944 10802 6008
rect 10819 5944 10883 6008
rect 10900 5944 10964 6008
rect 10981 5944 11045 6008
rect 11062 5944 11126 6008
rect 11143 5944 11207 6008
rect 11224 5944 11288 6008
rect 11305 5944 11369 6008
rect 11386 5944 11450 6008
rect 11467 5944 11531 6008
rect 11548 5944 11612 6008
rect 11629 5944 11693 6008
rect 11710 5944 11774 6008
rect 11791 5944 11855 6008
rect 11872 5944 11936 6008
rect 11953 5944 12017 6008
rect 12034 5944 12098 6008
rect 12115 5944 12179 6008
rect 12196 5944 12260 6008
rect 12277 5944 12341 6008
rect 12358 5944 12422 6008
rect 12439 5944 12503 6008
rect 12520 5944 12584 6008
rect 12601 5944 12665 6008
rect 12682 5944 12746 6008
rect 12763 5944 12827 6008
rect 12844 5944 12908 6008
rect 12925 5944 12989 6008
rect 13006 5944 13070 6008
rect 13087 5944 13151 6008
rect 13168 5944 13232 6008
rect 13249 5944 13313 6008
rect 13330 5944 13394 6008
rect 13411 5944 13475 6008
rect 13492 5944 13556 6008
rect 13573 5944 13637 6008
rect 13654 5944 13718 6008
rect 13735 5944 13799 6008
rect 13816 5944 13880 6008
rect 13897 5944 13961 6008
rect 13978 5944 14042 6008
rect 14059 5944 14123 6008
rect 14140 5944 14204 6008
rect 14221 5944 14285 6008
rect 14302 5944 14366 6008
rect 14383 5944 14447 6008
rect 14464 5944 14528 6008
rect 14545 5944 14609 6008
rect 14626 5944 14690 6008
rect 14707 5944 14771 6008
rect 14788 5944 14852 6008
rect 10084 5858 10148 5922
rect 10166 5858 10230 5922
rect 10248 5858 10312 5922
rect 10330 5858 10394 5922
rect 10412 5858 10476 5922
rect 10494 5858 10558 5922
rect 10576 5858 10640 5922
rect 10657 5858 10721 5922
rect 10738 5858 10802 5922
rect 10819 5858 10883 5922
rect 10900 5858 10964 5922
rect 10981 5858 11045 5922
rect 11062 5858 11126 5922
rect 11143 5858 11207 5922
rect 11224 5858 11288 5922
rect 11305 5858 11369 5922
rect 11386 5858 11450 5922
rect 11467 5858 11531 5922
rect 11548 5858 11612 5922
rect 11629 5858 11693 5922
rect 11710 5858 11774 5922
rect 11791 5858 11855 5922
rect 11872 5858 11936 5922
rect 11953 5858 12017 5922
rect 12034 5858 12098 5922
rect 12115 5858 12179 5922
rect 12196 5858 12260 5922
rect 12277 5858 12341 5922
rect 12358 5858 12422 5922
rect 12439 5858 12503 5922
rect 12520 5858 12584 5922
rect 12601 5858 12665 5922
rect 12682 5858 12746 5922
rect 12763 5858 12827 5922
rect 12844 5858 12908 5922
rect 12925 5858 12989 5922
rect 13006 5858 13070 5922
rect 13087 5858 13151 5922
rect 13168 5858 13232 5922
rect 13249 5858 13313 5922
rect 13330 5858 13394 5922
rect 13411 5858 13475 5922
rect 13492 5858 13556 5922
rect 13573 5858 13637 5922
rect 13654 5858 13718 5922
rect 13735 5858 13799 5922
rect 13816 5858 13880 5922
rect 13897 5858 13961 5922
rect 13978 5858 14042 5922
rect 14059 5858 14123 5922
rect 14140 5858 14204 5922
rect 14221 5858 14285 5922
rect 14302 5858 14366 5922
rect 14383 5858 14447 5922
rect 14464 5858 14528 5922
rect 14545 5858 14609 5922
rect 14626 5858 14690 5922
rect 14707 5858 14771 5922
rect 14788 5858 14852 5922
rect 10084 5772 10148 5836
rect 10166 5772 10230 5836
rect 10248 5772 10312 5836
rect 10330 5772 10394 5836
rect 10412 5772 10476 5836
rect 10494 5772 10558 5836
rect 10576 5772 10640 5836
rect 10657 5772 10721 5836
rect 10738 5772 10802 5836
rect 10819 5772 10883 5836
rect 10900 5772 10964 5836
rect 10981 5772 11045 5836
rect 11062 5772 11126 5836
rect 11143 5772 11207 5836
rect 11224 5772 11288 5836
rect 11305 5772 11369 5836
rect 11386 5772 11450 5836
rect 11467 5772 11531 5836
rect 11548 5772 11612 5836
rect 11629 5772 11693 5836
rect 11710 5772 11774 5836
rect 11791 5772 11855 5836
rect 11872 5772 11936 5836
rect 11953 5772 12017 5836
rect 12034 5772 12098 5836
rect 12115 5772 12179 5836
rect 12196 5772 12260 5836
rect 12277 5772 12341 5836
rect 12358 5772 12422 5836
rect 12439 5772 12503 5836
rect 12520 5772 12584 5836
rect 12601 5772 12665 5836
rect 12682 5772 12746 5836
rect 12763 5772 12827 5836
rect 12844 5772 12908 5836
rect 12925 5772 12989 5836
rect 13006 5772 13070 5836
rect 13087 5772 13151 5836
rect 13168 5772 13232 5836
rect 13249 5772 13313 5836
rect 13330 5772 13394 5836
rect 13411 5772 13475 5836
rect 13492 5772 13556 5836
rect 13573 5772 13637 5836
rect 13654 5772 13718 5836
rect 13735 5772 13799 5836
rect 13816 5772 13880 5836
rect 13897 5772 13961 5836
rect 13978 5772 14042 5836
rect 14059 5772 14123 5836
rect 14140 5772 14204 5836
rect 14221 5772 14285 5836
rect 14302 5772 14366 5836
rect 14383 5772 14447 5836
rect 14464 5772 14528 5836
rect 14545 5772 14609 5836
rect 14626 5772 14690 5836
rect 14707 5772 14771 5836
rect 14788 5772 14852 5836
rect 10084 5686 10148 5750
rect 10166 5686 10230 5750
rect 10248 5686 10312 5750
rect 10330 5686 10394 5750
rect 10412 5686 10476 5750
rect 10494 5686 10558 5750
rect 10576 5686 10640 5750
rect 10657 5686 10721 5750
rect 10738 5686 10802 5750
rect 10819 5686 10883 5750
rect 10900 5686 10964 5750
rect 10981 5686 11045 5750
rect 11062 5686 11126 5750
rect 11143 5686 11207 5750
rect 11224 5686 11288 5750
rect 11305 5686 11369 5750
rect 11386 5686 11450 5750
rect 11467 5686 11531 5750
rect 11548 5686 11612 5750
rect 11629 5686 11693 5750
rect 11710 5686 11774 5750
rect 11791 5686 11855 5750
rect 11872 5686 11936 5750
rect 11953 5686 12017 5750
rect 12034 5686 12098 5750
rect 12115 5686 12179 5750
rect 12196 5686 12260 5750
rect 12277 5686 12341 5750
rect 12358 5686 12422 5750
rect 12439 5686 12503 5750
rect 12520 5686 12584 5750
rect 12601 5686 12665 5750
rect 12682 5686 12746 5750
rect 12763 5686 12827 5750
rect 12844 5686 12908 5750
rect 12925 5686 12989 5750
rect 13006 5686 13070 5750
rect 13087 5686 13151 5750
rect 13168 5686 13232 5750
rect 13249 5686 13313 5750
rect 13330 5686 13394 5750
rect 13411 5686 13475 5750
rect 13492 5686 13556 5750
rect 13573 5686 13637 5750
rect 13654 5686 13718 5750
rect 13735 5686 13799 5750
rect 13816 5686 13880 5750
rect 13897 5686 13961 5750
rect 13978 5686 14042 5750
rect 14059 5686 14123 5750
rect 14140 5686 14204 5750
rect 14221 5686 14285 5750
rect 14302 5686 14366 5750
rect 14383 5686 14447 5750
rect 14464 5686 14528 5750
rect 14545 5686 14609 5750
rect 14626 5686 14690 5750
rect 14707 5686 14771 5750
rect 14788 5686 14852 5750
rect 10084 5600 10148 5664
rect 10166 5600 10230 5664
rect 10248 5600 10312 5664
rect 10330 5600 10394 5664
rect 10412 5600 10476 5664
rect 10494 5600 10558 5664
rect 10576 5600 10640 5664
rect 10657 5600 10721 5664
rect 10738 5600 10802 5664
rect 10819 5600 10883 5664
rect 10900 5600 10964 5664
rect 10981 5600 11045 5664
rect 11062 5600 11126 5664
rect 11143 5600 11207 5664
rect 11224 5600 11288 5664
rect 11305 5600 11369 5664
rect 11386 5600 11450 5664
rect 11467 5600 11531 5664
rect 11548 5600 11612 5664
rect 11629 5600 11693 5664
rect 11710 5600 11774 5664
rect 11791 5600 11855 5664
rect 11872 5600 11936 5664
rect 11953 5600 12017 5664
rect 12034 5600 12098 5664
rect 12115 5600 12179 5664
rect 12196 5600 12260 5664
rect 12277 5600 12341 5664
rect 12358 5600 12422 5664
rect 12439 5600 12503 5664
rect 12520 5600 12584 5664
rect 12601 5600 12665 5664
rect 12682 5600 12746 5664
rect 12763 5600 12827 5664
rect 12844 5600 12908 5664
rect 12925 5600 12989 5664
rect 13006 5600 13070 5664
rect 13087 5600 13151 5664
rect 13168 5600 13232 5664
rect 13249 5600 13313 5664
rect 13330 5600 13394 5664
rect 13411 5600 13475 5664
rect 13492 5600 13556 5664
rect 13573 5600 13637 5664
rect 13654 5600 13718 5664
rect 13735 5600 13799 5664
rect 13816 5600 13880 5664
rect 13897 5600 13961 5664
rect 13978 5600 14042 5664
rect 14059 5600 14123 5664
rect 14140 5600 14204 5664
rect 14221 5600 14285 5664
rect 14302 5600 14366 5664
rect 14383 5600 14447 5664
rect 14464 5600 14528 5664
rect 14545 5600 14609 5664
rect 14626 5600 14690 5664
rect 14707 5600 14771 5664
rect 14788 5600 14852 5664
rect 10084 5514 10148 5578
rect 10166 5514 10230 5578
rect 10248 5514 10312 5578
rect 10330 5514 10394 5578
rect 10412 5514 10476 5578
rect 10494 5514 10558 5578
rect 10576 5514 10640 5578
rect 10657 5514 10721 5578
rect 10738 5514 10802 5578
rect 10819 5514 10883 5578
rect 10900 5514 10964 5578
rect 10981 5514 11045 5578
rect 11062 5514 11126 5578
rect 11143 5514 11207 5578
rect 11224 5514 11288 5578
rect 11305 5514 11369 5578
rect 11386 5514 11450 5578
rect 11467 5514 11531 5578
rect 11548 5514 11612 5578
rect 11629 5514 11693 5578
rect 11710 5514 11774 5578
rect 11791 5514 11855 5578
rect 11872 5514 11936 5578
rect 11953 5514 12017 5578
rect 12034 5514 12098 5578
rect 12115 5514 12179 5578
rect 12196 5514 12260 5578
rect 12277 5514 12341 5578
rect 12358 5514 12422 5578
rect 12439 5514 12503 5578
rect 12520 5514 12584 5578
rect 12601 5514 12665 5578
rect 12682 5514 12746 5578
rect 12763 5514 12827 5578
rect 12844 5514 12908 5578
rect 12925 5514 12989 5578
rect 13006 5514 13070 5578
rect 13087 5514 13151 5578
rect 13168 5514 13232 5578
rect 13249 5514 13313 5578
rect 13330 5514 13394 5578
rect 13411 5514 13475 5578
rect 13492 5514 13556 5578
rect 13573 5514 13637 5578
rect 13654 5514 13718 5578
rect 13735 5514 13799 5578
rect 13816 5514 13880 5578
rect 13897 5514 13961 5578
rect 13978 5514 14042 5578
rect 14059 5514 14123 5578
rect 14140 5514 14204 5578
rect 14221 5514 14285 5578
rect 14302 5514 14366 5578
rect 14383 5514 14447 5578
rect 14464 5514 14528 5578
rect 14545 5514 14609 5578
rect 14626 5514 14690 5578
rect 14707 5514 14771 5578
rect 14788 5514 14852 5578
rect 10084 5428 10148 5492
rect 10166 5428 10230 5492
rect 10248 5428 10312 5492
rect 10330 5428 10394 5492
rect 10412 5428 10476 5492
rect 10494 5428 10558 5492
rect 10576 5428 10640 5492
rect 10657 5428 10721 5492
rect 10738 5428 10802 5492
rect 10819 5428 10883 5492
rect 10900 5428 10964 5492
rect 10981 5428 11045 5492
rect 11062 5428 11126 5492
rect 11143 5428 11207 5492
rect 11224 5428 11288 5492
rect 11305 5428 11369 5492
rect 11386 5428 11450 5492
rect 11467 5428 11531 5492
rect 11548 5428 11612 5492
rect 11629 5428 11693 5492
rect 11710 5428 11774 5492
rect 11791 5428 11855 5492
rect 11872 5428 11936 5492
rect 11953 5428 12017 5492
rect 12034 5428 12098 5492
rect 12115 5428 12179 5492
rect 12196 5428 12260 5492
rect 12277 5428 12341 5492
rect 12358 5428 12422 5492
rect 12439 5428 12503 5492
rect 12520 5428 12584 5492
rect 12601 5428 12665 5492
rect 12682 5428 12746 5492
rect 12763 5428 12827 5492
rect 12844 5428 12908 5492
rect 12925 5428 12989 5492
rect 13006 5428 13070 5492
rect 13087 5428 13151 5492
rect 13168 5428 13232 5492
rect 13249 5428 13313 5492
rect 13330 5428 13394 5492
rect 13411 5428 13475 5492
rect 13492 5428 13556 5492
rect 13573 5428 13637 5492
rect 13654 5428 13718 5492
rect 13735 5428 13799 5492
rect 13816 5428 13880 5492
rect 13897 5428 13961 5492
rect 13978 5428 14042 5492
rect 14059 5428 14123 5492
rect 14140 5428 14204 5492
rect 14221 5428 14285 5492
rect 14302 5428 14366 5492
rect 14383 5428 14447 5492
rect 14464 5428 14528 5492
rect 14545 5428 14609 5492
rect 14626 5428 14690 5492
rect 14707 5428 14771 5492
rect 14788 5428 14852 5492
rect 10084 5342 10148 5406
rect 10166 5342 10230 5406
rect 10248 5342 10312 5406
rect 10330 5342 10394 5406
rect 10412 5342 10476 5406
rect 10494 5342 10558 5406
rect 10576 5342 10640 5406
rect 10657 5342 10721 5406
rect 10738 5342 10802 5406
rect 10819 5342 10883 5406
rect 10900 5342 10964 5406
rect 10981 5342 11045 5406
rect 11062 5342 11126 5406
rect 11143 5342 11207 5406
rect 11224 5342 11288 5406
rect 11305 5342 11369 5406
rect 11386 5342 11450 5406
rect 11467 5342 11531 5406
rect 11548 5342 11612 5406
rect 11629 5342 11693 5406
rect 11710 5342 11774 5406
rect 11791 5342 11855 5406
rect 11872 5342 11936 5406
rect 11953 5342 12017 5406
rect 12034 5342 12098 5406
rect 12115 5342 12179 5406
rect 12196 5342 12260 5406
rect 12277 5342 12341 5406
rect 12358 5342 12422 5406
rect 12439 5342 12503 5406
rect 12520 5342 12584 5406
rect 12601 5342 12665 5406
rect 12682 5342 12746 5406
rect 12763 5342 12827 5406
rect 12844 5342 12908 5406
rect 12925 5342 12989 5406
rect 13006 5342 13070 5406
rect 13087 5342 13151 5406
rect 13168 5342 13232 5406
rect 13249 5342 13313 5406
rect 13330 5342 13394 5406
rect 13411 5342 13475 5406
rect 13492 5342 13556 5406
rect 13573 5342 13637 5406
rect 13654 5342 13718 5406
rect 13735 5342 13799 5406
rect 13816 5342 13880 5406
rect 13897 5342 13961 5406
rect 13978 5342 14042 5406
rect 14059 5342 14123 5406
rect 14140 5342 14204 5406
rect 14221 5342 14285 5406
rect 14302 5342 14366 5406
rect 14383 5342 14447 5406
rect 14464 5342 14528 5406
rect 14545 5342 14609 5406
rect 14626 5342 14690 5406
rect 14707 5342 14771 5406
rect 14788 5342 14852 5406
rect 10084 5256 10148 5320
rect 10166 5256 10230 5320
rect 10248 5256 10312 5320
rect 10330 5256 10394 5320
rect 10412 5256 10476 5320
rect 10494 5256 10558 5320
rect 10576 5256 10640 5320
rect 10657 5256 10721 5320
rect 10738 5256 10802 5320
rect 10819 5256 10883 5320
rect 10900 5256 10964 5320
rect 10981 5256 11045 5320
rect 11062 5256 11126 5320
rect 11143 5256 11207 5320
rect 11224 5256 11288 5320
rect 11305 5256 11369 5320
rect 11386 5256 11450 5320
rect 11467 5256 11531 5320
rect 11548 5256 11612 5320
rect 11629 5256 11693 5320
rect 11710 5256 11774 5320
rect 11791 5256 11855 5320
rect 11872 5256 11936 5320
rect 11953 5256 12017 5320
rect 12034 5256 12098 5320
rect 12115 5256 12179 5320
rect 12196 5256 12260 5320
rect 12277 5256 12341 5320
rect 12358 5256 12422 5320
rect 12439 5256 12503 5320
rect 12520 5256 12584 5320
rect 12601 5256 12665 5320
rect 12682 5256 12746 5320
rect 12763 5256 12827 5320
rect 12844 5256 12908 5320
rect 12925 5256 12989 5320
rect 13006 5256 13070 5320
rect 13087 5256 13151 5320
rect 13168 5256 13232 5320
rect 13249 5256 13313 5320
rect 13330 5256 13394 5320
rect 13411 5256 13475 5320
rect 13492 5256 13556 5320
rect 13573 5256 13637 5320
rect 13654 5256 13718 5320
rect 13735 5256 13799 5320
rect 13816 5256 13880 5320
rect 13897 5256 13961 5320
rect 13978 5256 14042 5320
rect 14059 5256 14123 5320
rect 14140 5256 14204 5320
rect 14221 5256 14285 5320
rect 14302 5256 14366 5320
rect 14383 5256 14447 5320
rect 14464 5256 14528 5320
rect 14545 5256 14609 5320
rect 14626 5256 14690 5320
rect 14707 5256 14771 5320
rect 14788 5256 14852 5320
rect 10084 5170 10148 5234
rect 10166 5170 10230 5234
rect 10248 5170 10312 5234
rect 10330 5170 10394 5234
rect 10412 5170 10476 5234
rect 10494 5170 10558 5234
rect 10576 5170 10640 5234
rect 10657 5170 10721 5234
rect 10738 5170 10802 5234
rect 10819 5170 10883 5234
rect 10900 5170 10964 5234
rect 10981 5170 11045 5234
rect 11062 5170 11126 5234
rect 11143 5170 11207 5234
rect 11224 5170 11288 5234
rect 11305 5170 11369 5234
rect 11386 5170 11450 5234
rect 11467 5170 11531 5234
rect 11548 5170 11612 5234
rect 11629 5170 11693 5234
rect 11710 5170 11774 5234
rect 11791 5170 11855 5234
rect 11872 5170 11936 5234
rect 11953 5170 12017 5234
rect 12034 5170 12098 5234
rect 12115 5170 12179 5234
rect 12196 5170 12260 5234
rect 12277 5170 12341 5234
rect 12358 5170 12422 5234
rect 12439 5170 12503 5234
rect 12520 5170 12584 5234
rect 12601 5170 12665 5234
rect 12682 5170 12746 5234
rect 12763 5170 12827 5234
rect 12844 5170 12908 5234
rect 12925 5170 12989 5234
rect 13006 5170 13070 5234
rect 13087 5170 13151 5234
rect 13168 5170 13232 5234
rect 13249 5170 13313 5234
rect 13330 5170 13394 5234
rect 13411 5170 13475 5234
rect 13492 5170 13556 5234
rect 13573 5170 13637 5234
rect 13654 5170 13718 5234
rect 13735 5170 13799 5234
rect 13816 5170 13880 5234
rect 13897 5170 13961 5234
rect 13978 5170 14042 5234
rect 14059 5170 14123 5234
rect 14140 5170 14204 5234
rect 14221 5170 14285 5234
rect 14302 5170 14366 5234
rect 14383 5170 14447 5234
rect 14464 5170 14528 5234
rect 14545 5170 14609 5234
rect 14626 5170 14690 5234
rect 14707 5170 14771 5234
rect 14788 5170 14852 5234
<< metal4 >>
rect 0 39984 254 40000
rect 0 39983 2695 39984
rect 0 39919 125 39983
rect 189 39919 205 39983
rect 269 39919 285 39983
rect 349 39919 365 39983
rect 429 39919 445 39983
rect 509 39919 525 39983
rect 589 39919 605 39983
rect 669 39919 685 39983
rect 749 39919 765 39983
rect 829 39919 845 39983
rect 909 39919 925 39983
rect 989 39919 1005 39983
rect 1069 39919 1085 39983
rect 1149 39919 1165 39983
rect 1229 39919 1245 39983
rect 1309 39919 1325 39983
rect 1389 39919 1405 39983
rect 1469 39919 1485 39983
rect 1549 39919 1565 39983
rect 1629 39919 1645 39983
rect 1709 39919 1725 39983
rect 1789 39919 1805 39983
rect 1869 39919 1885 39983
rect 1949 39919 1965 39983
rect 2029 39919 2045 39983
rect 2109 39919 2125 39983
rect 2189 39919 2205 39983
rect 2269 39919 2285 39983
rect 2349 39919 2365 39983
rect 2429 39919 2445 39983
rect 2509 39919 2525 39983
rect 2589 39919 2605 39983
rect 2669 39919 2695 39983
rect 0 39902 2695 39919
rect 0 39838 125 39902
rect 189 39838 205 39902
rect 269 39838 285 39902
rect 349 39838 365 39902
rect 429 39838 445 39902
rect 509 39838 525 39902
rect 589 39838 605 39902
rect 669 39838 685 39902
rect 749 39838 765 39902
rect 829 39838 845 39902
rect 909 39838 925 39902
rect 989 39838 1005 39902
rect 1069 39838 1085 39902
rect 1149 39838 1165 39902
rect 1229 39838 1245 39902
rect 1309 39838 1325 39902
rect 1389 39838 1405 39902
rect 1469 39838 1485 39902
rect 1549 39838 1565 39902
rect 1629 39838 1645 39902
rect 1709 39838 1725 39902
rect 1789 39838 1805 39902
rect 1869 39838 1885 39902
rect 1949 39838 1965 39902
rect 2029 39838 2045 39902
rect 2109 39838 2125 39902
rect 2189 39838 2205 39902
rect 2269 39838 2285 39902
rect 2349 39838 2365 39902
rect 2429 39838 2445 39902
rect 2509 39838 2525 39902
rect 2589 39838 2605 39902
rect 2669 39838 2695 39902
rect 0 39821 2695 39838
rect 0 39757 125 39821
rect 189 39757 205 39821
rect 269 39757 285 39821
rect 349 39757 365 39821
rect 429 39757 445 39821
rect 509 39757 525 39821
rect 589 39757 605 39821
rect 669 39757 685 39821
rect 749 39757 765 39821
rect 829 39757 845 39821
rect 909 39757 925 39821
rect 989 39757 1005 39821
rect 1069 39757 1085 39821
rect 1149 39757 1165 39821
rect 1229 39757 1245 39821
rect 1309 39757 1325 39821
rect 1389 39757 1405 39821
rect 1469 39757 1485 39821
rect 1549 39757 1565 39821
rect 1629 39757 1645 39821
rect 1709 39757 1725 39821
rect 1789 39757 1805 39821
rect 1869 39757 1885 39821
rect 1949 39757 1965 39821
rect 2029 39757 2045 39821
rect 2109 39757 2125 39821
rect 2189 39757 2205 39821
rect 2269 39757 2285 39821
rect 2349 39757 2365 39821
rect 2429 39757 2445 39821
rect 2509 39757 2525 39821
rect 2589 39757 2605 39821
rect 2669 39757 2695 39821
rect 0 39740 2695 39757
rect 0 39676 125 39740
rect 189 39676 205 39740
rect 269 39676 285 39740
rect 349 39676 365 39740
rect 429 39676 445 39740
rect 509 39676 525 39740
rect 589 39676 605 39740
rect 669 39676 685 39740
rect 749 39676 765 39740
rect 829 39676 845 39740
rect 909 39676 925 39740
rect 989 39676 1005 39740
rect 1069 39676 1085 39740
rect 1149 39676 1165 39740
rect 1229 39676 1245 39740
rect 1309 39676 1325 39740
rect 1389 39676 1405 39740
rect 1469 39676 1485 39740
rect 1549 39676 1565 39740
rect 1629 39676 1645 39740
rect 1709 39676 1725 39740
rect 1789 39676 1805 39740
rect 1869 39676 1885 39740
rect 1949 39676 1965 39740
rect 2029 39676 2045 39740
rect 2109 39676 2125 39740
rect 2189 39676 2205 39740
rect 2269 39676 2285 39740
rect 2349 39676 2365 39740
rect 2429 39676 2445 39740
rect 2509 39676 2525 39740
rect 2589 39676 2605 39740
rect 2669 39676 2695 39740
rect 0 39659 2695 39676
rect 0 39595 125 39659
rect 189 39595 205 39659
rect 269 39595 285 39659
rect 349 39595 365 39659
rect 429 39595 445 39659
rect 509 39595 525 39659
rect 589 39595 605 39659
rect 669 39595 685 39659
rect 749 39595 765 39659
rect 829 39595 845 39659
rect 909 39595 925 39659
rect 989 39595 1005 39659
rect 1069 39595 1085 39659
rect 1149 39595 1165 39659
rect 1229 39595 1245 39659
rect 1309 39595 1325 39659
rect 1389 39595 1405 39659
rect 1469 39595 1485 39659
rect 1549 39595 1565 39659
rect 1629 39595 1645 39659
rect 1709 39595 1725 39659
rect 1789 39595 1805 39659
rect 1869 39595 1885 39659
rect 1949 39595 1965 39659
rect 2029 39595 2045 39659
rect 2109 39595 2125 39659
rect 2189 39595 2205 39659
rect 2269 39595 2285 39659
rect 2349 39595 2365 39659
rect 2429 39595 2445 39659
rect 2509 39595 2525 39659
rect 2589 39595 2605 39659
rect 2669 39595 2695 39659
rect 0 39578 2695 39595
rect 0 39514 125 39578
rect 189 39514 205 39578
rect 269 39514 285 39578
rect 349 39514 365 39578
rect 429 39514 445 39578
rect 509 39514 525 39578
rect 589 39514 605 39578
rect 669 39514 685 39578
rect 749 39514 765 39578
rect 829 39514 845 39578
rect 909 39514 925 39578
rect 989 39514 1005 39578
rect 1069 39514 1085 39578
rect 1149 39514 1165 39578
rect 1229 39514 1245 39578
rect 1309 39514 1325 39578
rect 1389 39514 1405 39578
rect 1469 39514 1485 39578
rect 1549 39514 1565 39578
rect 1629 39514 1645 39578
rect 1709 39514 1725 39578
rect 1789 39514 1805 39578
rect 1869 39514 1885 39578
rect 1949 39514 1965 39578
rect 2029 39514 2045 39578
rect 2109 39514 2125 39578
rect 2189 39514 2205 39578
rect 2269 39514 2285 39578
rect 2349 39514 2365 39578
rect 2429 39514 2445 39578
rect 2509 39514 2525 39578
rect 2589 39514 2605 39578
rect 2669 39514 2695 39578
rect 0 39497 2695 39514
rect 0 39433 125 39497
rect 189 39433 205 39497
rect 269 39433 285 39497
rect 349 39433 365 39497
rect 429 39433 445 39497
rect 509 39433 525 39497
rect 589 39433 605 39497
rect 669 39433 685 39497
rect 749 39433 765 39497
rect 829 39433 845 39497
rect 909 39433 925 39497
rect 989 39433 1005 39497
rect 1069 39433 1085 39497
rect 1149 39433 1165 39497
rect 1229 39433 1245 39497
rect 1309 39433 1325 39497
rect 1389 39433 1405 39497
rect 1469 39433 1485 39497
rect 1549 39433 1565 39497
rect 1629 39433 1645 39497
rect 1709 39433 1725 39497
rect 1789 39433 1805 39497
rect 1869 39433 1885 39497
rect 1949 39433 1965 39497
rect 2029 39433 2045 39497
rect 2109 39433 2125 39497
rect 2189 39433 2205 39497
rect 2269 39433 2285 39497
rect 2349 39433 2365 39497
rect 2429 39433 2445 39497
rect 2509 39433 2525 39497
rect 2589 39433 2605 39497
rect 2669 39433 2695 39497
rect 2726 39982 12265 39986
rect 14746 39984 15000 40000
rect 2726 39918 2727 39982
rect 2791 39918 2808 39982
rect 2872 39918 2889 39982
rect 2953 39918 2970 39982
rect 3034 39918 3051 39982
rect 3115 39918 3132 39982
rect 3196 39918 3213 39982
rect 3277 39918 3294 39982
rect 3358 39918 3375 39982
rect 3439 39918 3456 39982
rect 3520 39918 3537 39982
rect 3601 39918 3618 39982
rect 3682 39918 3699 39982
rect 3763 39918 3780 39982
rect 3844 39918 3861 39982
rect 3925 39918 3942 39982
rect 4006 39918 4023 39982
rect 4087 39918 4104 39982
rect 4168 39918 4185 39982
rect 4249 39918 4266 39982
rect 4330 39918 4347 39982
rect 4411 39918 4428 39982
rect 4492 39918 4509 39982
rect 4573 39918 4590 39982
rect 4654 39918 4671 39982
rect 4735 39918 4752 39982
rect 4816 39918 4833 39982
rect 4897 39918 4914 39982
rect 4978 39918 4995 39982
rect 5059 39918 5076 39982
rect 5140 39918 5157 39982
rect 5221 39918 5238 39982
rect 5302 39918 5319 39982
rect 5383 39918 5400 39982
rect 2726 39902 5400 39918
rect 2726 39838 2727 39902
rect 2791 39838 2808 39902
rect 2872 39838 2889 39902
rect 2953 39838 2970 39902
rect 3034 39838 3051 39902
rect 3115 39838 3132 39902
rect 3196 39838 3213 39902
rect 3277 39838 3294 39902
rect 3358 39838 3375 39902
rect 3439 39838 3456 39902
rect 3520 39838 3537 39902
rect 3601 39838 3618 39902
rect 3682 39838 3699 39902
rect 3763 39838 3780 39902
rect 3844 39838 3861 39902
rect 3925 39838 3942 39902
rect 4006 39838 4023 39902
rect 4087 39838 4104 39902
rect 4168 39838 4185 39902
rect 4249 39838 4266 39902
rect 4330 39838 4347 39902
rect 4411 39838 4428 39902
rect 4492 39838 4509 39902
rect 4573 39838 4590 39902
rect 4654 39838 4671 39902
rect 4735 39838 4752 39902
rect 4816 39838 4833 39902
rect 4897 39838 4914 39902
rect 4978 39838 4995 39902
rect 5059 39838 5076 39902
rect 5140 39838 5157 39902
rect 5221 39838 5238 39902
rect 5302 39838 5319 39902
rect 5383 39838 5400 39902
rect 2726 39822 5400 39838
rect 2726 39758 2727 39822
rect 2791 39758 2808 39822
rect 2872 39758 2889 39822
rect 2953 39758 2970 39822
rect 3034 39758 3051 39822
rect 3115 39758 3132 39822
rect 3196 39758 3213 39822
rect 3277 39758 3294 39822
rect 3358 39758 3375 39822
rect 3439 39758 3456 39822
rect 3520 39758 3537 39822
rect 3601 39758 3618 39822
rect 3682 39758 3699 39822
rect 3763 39758 3780 39822
rect 3844 39758 3861 39822
rect 3925 39758 3942 39822
rect 4006 39758 4023 39822
rect 4087 39758 4104 39822
rect 4168 39758 4185 39822
rect 4249 39758 4266 39822
rect 4330 39758 4347 39822
rect 4411 39758 4428 39822
rect 4492 39758 4509 39822
rect 4573 39758 4590 39822
rect 4654 39758 4671 39822
rect 4735 39758 4752 39822
rect 4816 39758 4833 39822
rect 4897 39758 4914 39822
rect 4978 39758 4995 39822
rect 5059 39758 5076 39822
rect 5140 39758 5157 39822
rect 5221 39758 5238 39822
rect 5302 39758 5319 39822
rect 5383 39758 5400 39822
rect 2726 39742 5400 39758
rect 2726 39678 2727 39742
rect 2791 39678 2808 39742
rect 2872 39678 2889 39742
rect 2953 39678 2970 39742
rect 3034 39678 3051 39742
rect 3115 39678 3132 39742
rect 3196 39678 3213 39742
rect 3277 39678 3294 39742
rect 3358 39678 3375 39742
rect 3439 39678 3456 39742
rect 3520 39678 3537 39742
rect 3601 39678 3618 39742
rect 3682 39678 3699 39742
rect 3763 39678 3780 39742
rect 3844 39678 3861 39742
rect 3925 39678 3942 39742
rect 4006 39678 4023 39742
rect 4087 39678 4104 39742
rect 4168 39678 4185 39742
rect 4249 39678 4266 39742
rect 4330 39678 4347 39742
rect 4411 39678 4428 39742
rect 4492 39678 4509 39742
rect 4573 39678 4590 39742
rect 4654 39678 4671 39742
rect 4735 39678 4752 39742
rect 4816 39678 4833 39742
rect 4897 39678 4914 39742
rect 4978 39678 4995 39742
rect 5059 39678 5076 39742
rect 5140 39678 5157 39742
rect 5221 39678 5238 39742
rect 5302 39678 5319 39742
rect 5383 39678 5400 39742
rect 2726 39662 5400 39678
rect 2726 39598 2727 39662
rect 2791 39598 2808 39662
rect 2872 39598 2889 39662
rect 2953 39598 2970 39662
rect 3034 39598 3051 39662
rect 3115 39598 3132 39662
rect 3196 39598 3213 39662
rect 3277 39598 3294 39662
rect 3358 39598 3375 39662
rect 3439 39598 3456 39662
rect 3520 39598 3537 39662
rect 3601 39598 3618 39662
rect 3682 39598 3699 39662
rect 3763 39598 3780 39662
rect 3844 39598 3861 39662
rect 3925 39598 3942 39662
rect 4006 39598 4023 39662
rect 4087 39598 4104 39662
rect 4168 39598 4185 39662
rect 4249 39598 4266 39662
rect 4330 39598 4347 39662
rect 4411 39598 4428 39662
rect 4492 39598 4509 39662
rect 4573 39598 4590 39662
rect 4654 39598 4671 39662
rect 4735 39598 4752 39662
rect 4816 39598 4833 39662
rect 4897 39598 4914 39662
rect 4978 39598 4995 39662
rect 5059 39598 5076 39662
rect 5140 39598 5157 39662
rect 5221 39598 5238 39662
rect 5302 39598 5319 39662
rect 5383 39598 5400 39662
rect 2726 39582 5400 39598
rect 2726 39518 2727 39582
rect 2791 39518 2808 39582
rect 2872 39518 2889 39582
rect 2953 39518 2970 39582
rect 3034 39518 3051 39582
rect 3115 39518 3132 39582
rect 3196 39518 3213 39582
rect 3277 39518 3294 39582
rect 3358 39518 3375 39582
rect 3439 39518 3456 39582
rect 3520 39518 3537 39582
rect 3601 39518 3618 39582
rect 3682 39518 3699 39582
rect 3763 39518 3780 39582
rect 3844 39518 3861 39582
rect 3925 39518 3942 39582
rect 4006 39518 4023 39582
rect 4087 39518 4104 39582
rect 4168 39518 4185 39582
rect 4249 39518 4266 39582
rect 4330 39518 4347 39582
rect 4411 39518 4428 39582
rect 4492 39518 4509 39582
rect 4573 39518 4590 39582
rect 4654 39518 4671 39582
rect 4735 39518 4752 39582
rect 4816 39518 4833 39582
rect 4897 39518 4914 39582
rect 4978 39518 4995 39582
rect 5059 39518 5076 39582
rect 5140 39518 5157 39582
rect 5221 39518 5238 39582
rect 5302 39518 5319 39582
rect 5383 39518 5400 39582
rect 2726 39502 5400 39518
rect 2726 39438 2727 39502
rect 2791 39438 2808 39502
rect 2872 39438 2889 39502
rect 2953 39438 2970 39502
rect 3034 39438 3051 39502
rect 3115 39438 3132 39502
rect 3196 39438 3213 39502
rect 3277 39438 3294 39502
rect 3358 39438 3375 39502
rect 3439 39438 3456 39502
rect 3520 39438 3537 39502
rect 3601 39438 3618 39502
rect 3682 39438 3699 39502
rect 3763 39438 3780 39502
rect 3844 39438 3861 39502
rect 3925 39438 3942 39502
rect 4006 39438 4023 39502
rect 4087 39438 4104 39502
rect 4168 39438 4185 39502
rect 4249 39438 4266 39502
rect 4330 39438 4347 39502
rect 4411 39438 4428 39502
rect 4492 39438 4509 39502
rect 4573 39438 4590 39502
rect 4654 39438 4671 39502
rect 4735 39438 4752 39502
rect 4816 39438 4833 39502
rect 4897 39438 4914 39502
rect 4978 39438 4995 39502
rect 5059 39438 5076 39502
rect 5140 39438 5157 39502
rect 5221 39438 5238 39502
rect 5302 39438 5319 39502
rect 5383 39438 5400 39502
rect 12264 39438 12265 39982
rect 2726 39434 12265 39438
rect 12301 39983 15000 39984
rect 12301 39919 12306 39983
rect 12370 39919 12386 39983
rect 12450 39919 12466 39983
rect 12530 39919 12546 39983
rect 12610 39919 12626 39983
rect 12690 39919 12706 39983
rect 12770 39919 12786 39983
rect 12850 39919 12866 39983
rect 12930 39919 12946 39983
rect 13010 39919 13026 39983
rect 13090 39919 13106 39983
rect 13170 39919 13186 39983
rect 13250 39919 13266 39983
rect 13330 39919 13346 39983
rect 13410 39919 13426 39983
rect 13490 39919 13506 39983
rect 13570 39919 13586 39983
rect 13650 39919 13666 39983
rect 13730 39919 13746 39983
rect 13810 39919 13826 39983
rect 13890 39919 13906 39983
rect 13970 39919 13986 39983
rect 14050 39919 14066 39983
rect 14130 39919 14146 39983
rect 14210 39919 14226 39983
rect 14290 39919 14306 39983
rect 14370 39919 14386 39983
rect 14450 39919 14466 39983
rect 14530 39919 14546 39983
rect 14610 39919 14626 39983
rect 14690 39919 14706 39983
rect 14770 39919 14786 39983
rect 14850 39919 15000 39983
rect 12301 39902 15000 39919
rect 12301 39838 12306 39902
rect 12370 39838 12386 39902
rect 12450 39838 12466 39902
rect 12530 39838 12546 39902
rect 12610 39838 12626 39902
rect 12690 39838 12706 39902
rect 12770 39838 12786 39902
rect 12850 39838 12866 39902
rect 12930 39838 12946 39902
rect 13010 39838 13026 39902
rect 13090 39838 13106 39902
rect 13170 39838 13186 39902
rect 13250 39838 13266 39902
rect 13330 39838 13346 39902
rect 13410 39838 13426 39902
rect 13490 39838 13506 39902
rect 13570 39838 13586 39902
rect 13650 39838 13666 39902
rect 13730 39838 13746 39902
rect 13810 39838 13826 39902
rect 13890 39838 13906 39902
rect 13970 39838 13986 39902
rect 14050 39838 14066 39902
rect 14130 39838 14146 39902
rect 14210 39838 14226 39902
rect 14290 39838 14306 39902
rect 14370 39838 14386 39902
rect 14450 39838 14466 39902
rect 14530 39838 14546 39902
rect 14610 39838 14626 39902
rect 14690 39838 14706 39902
rect 14770 39838 14786 39902
rect 14850 39838 15000 39902
rect 12301 39821 15000 39838
rect 12301 39757 12306 39821
rect 12370 39757 12386 39821
rect 12450 39757 12466 39821
rect 12530 39757 12546 39821
rect 12610 39757 12626 39821
rect 12690 39757 12706 39821
rect 12770 39757 12786 39821
rect 12850 39757 12866 39821
rect 12930 39757 12946 39821
rect 13010 39757 13026 39821
rect 13090 39757 13106 39821
rect 13170 39757 13186 39821
rect 13250 39757 13266 39821
rect 13330 39757 13346 39821
rect 13410 39757 13426 39821
rect 13490 39757 13506 39821
rect 13570 39757 13586 39821
rect 13650 39757 13666 39821
rect 13730 39757 13746 39821
rect 13810 39757 13826 39821
rect 13890 39757 13906 39821
rect 13970 39757 13986 39821
rect 14050 39757 14066 39821
rect 14130 39757 14146 39821
rect 14210 39757 14226 39821
rect 14290 39757 14306 39821
rect 14370 39757 14386 39821
rect 14450 39757 14466 39821
rect 14530 39757 14546 39821
rect 14610 39757 14626 39821
rect 14690 39757 14706 39821
rect 14770 39757 14786 39821
rect 14850 39757 15000 39821
rect 12301 39740 15000 39757
rect 12301 39676 12306 39740
rect 12370 39676 12386 39740
rect 12450 39676 12466 39740
rect 12530 39676 12546 39740
rect 12610 39676 12626 39740
rect 12690 39676 12706 39740
rect 12770 39676 12786 39740
rect 12850 39676 12866 39740
rect 12930 39676 12946 39740
rect 13010 39676 13026 39740
rect 13090 39676 13106 39740
rect 13170 39676 13186 39740
rect 13250 39676 13266 39740
rect 13330 39676 13346 39740
rect 13410 39676 13426 39740
rect 13490 39676 13506 39740
rect 13570 39676 13586 39740
rect 13650 39676 13666 39740
rect 13730 39676 13746 39740
rect 13810 39676 13826 39740
rect 13890 39676 13906 39740
rect 13970 39676 13986 39740
rect 14050 39676 14066 39740
rect 14130 39676 14146 39740
rect 14210 39676 14226 39740
rect 14290 39676 14306 39740
rect 14370 39676 14386 39740
rect 14450 39676 14466 39740
rect 14530 39676 14546 39740
rect 14610 39676 14626 39740
rect 14690 39676 14706 39740
rect 14770 39676 14786 39740
rect 14850 39676 15000 39740
rect 12301 39659 15000 39676
rect 12301 39595 12306 39659
rect 12370 39595 12386 39659
rect 12450 39595 12466 39659
rect 12530 39595 12546 39659
rect 12610 39595 12626 39659
rect 12690 39595 12706 39659
rect 12770 39595 12786 39659
rect 12850 39595 12866 39659
rect 12930 39595 12946 39659
rect 13010 39595 13026 39659
rect 13090 39595 13106 39659
rect 13170 39595 13186 39659
rect 13250 39595 13266 39659
rect 13330 39595 13346 39659
rect 13410 39595 13426 39659
rect 13490 39595 13506 39659
rect 13570 39595 13586 39659
rect 13650 39595 13666 39659
rect 13730 39595 13746 39659
rect 13810 39595 13826 39659
rect 13890 39595 13906 39659
rect 13970 39595 13986 39659
rect 14050 39595 14066 39659
rect 14130 39595 14146 39659
rect 14210 39595 14226 39659
rect 14290 39595 14306 39659
rect 14370 39595 14386 39659
rect 14450 39595 14466 39659
rect 14530 39595 14546 39659
rect 14610 39595 14626 39659
rect 14690 39595 14706 39659
rect 14770 39595 14786 39659
rect 14850 39595 15000 39659
rect 12301 39578 15000 39595
rect 12301 39514 12306 39578
rect 12370 39514 12386 39578
rect 12450 39514 12466 39578
rect 12530 39514 12546 39578
rect 12610 39514 12626 39578
rect 12690 39514 12706 39578
rect 12770 39514 12786 39578
rect 12850 39514 12866 39578
rect 12930 39514 12946 39578
rect 13010 39514 13026 39578
rect 13090 39514 13106 39578
rect 13170 39514 13186 39578
rect 13250 39514 13266 39578
rect 13330 39514 13346 39578
rect 13410 39514 13426 39578
rect 13490 39514 13506 39578
rect 13570 39514 13586 39578
rect 13650 39514 13666 39578
rect 13730 39514 13746 39578
rect 13810 39514 13826 39578
rect 13890 39514 13906 39578
rect 13970 39514 13986 39578
rect 14050 39514 14066 39578
rect 14130 39514 14146 39578
rect 14210 39514 14226 39578
rect 14290 39514 14306 39578
rect 14370 39514 14386 39578
rect 14450 39514 14466 39578
rect 14530 39514 14546 39578
rect 14610 39514 14626 39578
rect 14690 39514 14706 39578
rect 14770 39514 14786 39578
rect 14850 39514 15000 39578
rect 12301 39497 15000 39514
rect 0 39416 2695 39433
rect 0 39352 125 39416
rect 189 39352 205 39416
rect 269 39352 285 39416
rect 349 39352 365 39416
rect 429 39352 445 39416
rect 509 39352 525 39416
rect 589 39352 605 39416
rect 669 39352 685 39416
rect 749 39352 765 39416
rect 829 39352 845 39416
rect 909 39352 925 39416
rect 989 39352 1005 39416
rect 1069 39352 1085 39416
rect 1149 39352 1165 39416
rect 1229 39352 1245 39416
rect 1309 39352 1325 39416
rect 1389 39352 1405 39416
rect 1469 39352 1485 39416
rect 1549 39352 1565 39416
rect 1629 39352 1645 39416
rect 1709 39352 1725 39416
rect 1789 39352 1805 39416
rect 1869 39352 1885 39416
rect 1949 39352 1965 39416
rect 2029 39352 2045 39416
rect 2109 39352 2125 39416
rect 2189 39352 2205 39416
rect 2269 39352 2285 39416
rect 2349 39352 2365 39416
rect 2429 39352 2445 39416
rect 2509 39352 2525 39416
rect 2589 39352 2605 39416
rect 2669 39352 2695 39416
rect 12301 39433 12306 39497
rect 12370 39433 12386 39497
rect 12450 39433 12466 39497
rect 12530 39433 12546 39497
rect 12610 39433 12626 39497
rect 12690 39433 12706 39497
rect 12770 39433 12786 39497
rect 12850 39433 12866 39497
rect 12930 39433 12946 39497
rect 13010 39433 13026 39497
rect 13090 39433 13106 39497
rect 13170 39433 13186 39497
rect 13250 39433 13266 39497
rect 13330 39433 13346 39497
rect 13410 39433 13426 39497
rect 13490 39433 13506 39497
rect 13570 39433 13586 39497
rect 13650 39433 13666 39497
rect 13730 39433 13746 39497
rect 13810 39433 13826 39497
rect 13890 39433 13906 39497
rect 13970 39433 13986 39497
rect 14050 39433 14066 39497
rect 14130 39433 14146 39497
rect 14210 39433 14226 39497
rect 14290 39433 14306 39497
rect 14370 39433 14386 39497
rect 14450 39433 14466 39497
rect 14530 39433 14546 39497
rect 14610 39433 14626 39497
rect 14690 39433 14706 39497
rect 14770 39433 14786 39497
rect 14850 39433 15000 39497
rect 12301 39416 15000 39433
rect 0 39335 2695 39352
rect 0 39271 125 39335
rect 189 39271 205 39335
rect 269 39271 285 39335
rect 349 39271 365 39335
rect 429 39271 445 39335
rect 509 39271 525 39335
rect 589 39271 605 39335
rect 669 39271 685 39335
rect 749 39271 765 39335
rect 829 39271 845 39335
rect 909 39271 925 39335
rect 989 39271 1005 39335
rect 1069 39271 1085 39335
rect 1149 39271 1165 39335
rect 1229 39271 1245 39335
rect 1309 39271 1325 39335
rect 1389 39271 1405 39335
rect 1469 39271 1485 39335
rect 1549 39271 1565 39335
rect 1629 39271 1645 39335
rect 1709 39271 1725 39335
rect 1789 39271 1805 39335
rect 1869 39271 1885 39335
rect 1949 39271 1965 39335
rect 2029 39271 2045 39335
rect 2109 39271 2125 39335
rect 2189 39271 2205 39335
rect 2269 39271 2285 39335
rect 2349 39271 2365 39335
rect 2429 39271 2445 39335
rect 2509 39271 2525 39335
rect 2589 39271 2605 39335
rect 2669 39271 2695 39335
rect 0 39254 2695 39271
rect 0 39190 125 39254
rect 189 39190 205 39254
rect 269 39190 285 39254
rect 349 39190 365 39254
rect 429 39190 445 39254
rect 509 39190 525 39254
rect 589 39190 605 39254
rect 669 39190 685 39254
rect 749 39190 765 39254
rect 829 39190 845 39254
rect 909 39190 925 39254
rect 989 39190 1005 39254
rect 1069 39190 1085 39254
rect 1149 39190 1165 39254
rect 1229 39190 1245 39254
rect 1309 39190 1325 39254
rect 1389 39190 1405 39254
rect 1469 39190 1485 39254
rect 1549 39190 1565 39254
rect 1629 39190 1645 39254
rect 1709 39190 1725 39254
rect 1789 39190 1805 39254
rect 1869 39190 1885 39254
rect 1949 39190 1965 39254
rect 2029 39190 2045 39254
rect 2109 39190 2125 39254
rect 2189 39190 2205 39254
rect 2269 39190 2285 39254
rect 2349 39190 2365 39254
rect 2429 39190 2445 39254
rect 2509 39190 2525 39254
rect 2589 39190 2605 39254
rect 2669 39190 2695 39254
rect 2719 39393 2851 39394
rect 2719 39329 2753 39393
rect 2817 39329 2851 39393
rect 2719 39311 2851 39329
rect 2719 39247 2753 39311
rect 2817 39247 2851 39311
rect 2719 39246 2851 39247
rect 12136 39393 12268 39394
rect 12136 39329 12170 39393
rect 12234 39329 12268 39393
rect 12136 39311 12268 39329
rect 12136 39247 12170 39311
rect 12234 39247 12268 39311
rect 12136 39246 12268 39247
rect 12301 39352 12306 39416
rect 12370 39352 12386 39416
rect 12450 39352 12466 39416
rect 12530 39352 12546 39416
rect 12610 39352 12626 39416
rect 12690 39352 12706 39416
rect 12770 39352 12786 39416
rect 12850 39352 12866 39416
rect 12930 39352 12946 39416
rect 13010 39352 13026 39416
rect 13090 39352 13106 39416
rect 13170 39352 13186 39416
rect 13250 39352 13266 39416
rect 13330 39352 13346 39416
rect 13410 39352 13426 39416
rect 13490 39352 13506 39416
rect 13570 39352 13586 39416
rect 13650 39352 13666 39416
rect 13730 39352 13746 39416
rect 13810 39352 13826 39416
rect 13890 39352 13906 39416
rect 13970 39352 13986 39416
rect 14050 39352 14066 39416
rect 14130 39352 14146 39416
rect 14210 39352 14226 39416
rect 14290 39352 14306 39416
rect 14370 39352 14386 39416
rect 14450 39352 14466 39416
rect 14530 39352 14546 39416
rect 14610 39352 14626 39416
rect 14690 39352 14706 39416
rect 14770 39352 14786 39416
rect 14850 39352 15000 39416
rect 12301 39335 15000 39352
rect 12301 39271 12306 39335
rect 12370 39271 12386 39335
rect 12450 39271 12466 39335
rect 12530 39271 12546 39335
rect 12610 39271 12626 39335
rect 12690 39271 12706 39335
rect 12770 39271 12786 39335
rect 12850 39271 12866 39335
rect 12930 39271 12946 39335
rect 13010 39271 13026 39335
rect 13090 39271 13106 39335
rect 13170 39271 13186 39335
rect 13250 39271 13266 39335
rect 13330 39271 13346 39335
rect 13410 39271 13426 39335
rect 13490 39271 13506 39335
rect 13570 39271 13586 39335
rect 13650 39271 13666 39335
rect 13730 39271 13746 39335
rect 13810 39271 13826 39335
rect 13890 39271 13906 39335
rect 13970 39271 13986 39335
rect 14050 39271 14066 39335
rect 14130 39271 14146 39335
rect 14210 39271 14226 39335
rect 14290 39271 14306 39335
rect 14370 39271 14386 39335
rect 14450 39271 14466 39335
rect 14530 39271 14546 39335
rect 14610 39271 14626 39335
rect 14690 39271 14706 39335
rect 14770 39271 14786 39335
rect 14850 39271 15000 39335
rect 12301 39254 15000 39271
rect 0 39173 2695 39190
rect 0 39109 125 39173
rect 189 39109 205 39173
rect 269 39109 285 39173
rect 349 39109 365 39173
rect 429 39109 445 39173
rect 509 39109 525 39173
rect 589 39109 605 39173
rect 669 39109 685 39173
rect 749 39109 765 39173
rect 829 39109 845 39173
rect 909 39109 925 39173
rect 989 39109 1005 39173
rect 1069 39109 1085 39173
rect 1149 39109 1165 39173
rect 1229 39109 1245 39173
rect 1309 39109 1325 39173
rect 1389 39109 1405 39173
rect 1469 39109 1485 39173
rect 1549 39109 1565 39173
rect 1629 39109 1645 39173
rect 1709 39109 1725 39173
rect 1789 39109 1805 39173
rect 1869 39109 1885 39173
rect 1949 39109 1965 39173
rect 2029 39109 2045 39173
rect 2109 39109 2125 39173
rect 2189 39109 2205 39173
rect 2269 39109 2285 39173
rect 2349 39109 2365 39173
rect 2429 39109 2445 39173
rect 2509 39109 2525 39173
rect 2589 39109 2605 39173
rect 2669 39109 2695 39173
rect 0 39092 2695 39109
rect 0 39028 125 39092
rect 189 39028 205 39092
rect 269 39028 285 39092
rect 349 39028 365 39092
rect 429 39028 445 39092
rect 509 39028 525 39092
rect 589 39028 605 39092
rect 669 39028 685 39092
rect 749 39028 765 39092
rect 829 39028 845 39092
rect 909 39028 925 39092
rect 989 39028 1005 39092
rect 1069 39028 1085 39092
rect 1149 39028 1165 39092
rect 1229 39028 1245 39092
rect 1309 39028 1325 39092
rect 1389 39028 1405 39092
rect 1469 39028 1485 39092
rect 1549 39028 1565 39092
rect 1629 39028 1645 39092
rect 1709 39028 1725 39092
rect 1789 39028 1805 39092
rect 1869 39028 1885 39092
rect 1949 39028 1965 39092
rect 2029 39028 2045 39092
rect 2109 39028 2125 39092
rect 2189 39028 2205 39092
rect 2269 39028 2285 39092
rect 2349 39028 2365 39092
rect 2429 39028 2445 39092
rect 2509 39028 2525 39092
rect 2589 39028 2605 39092
rect 2669 39028 2695 39092
rect 0 39011 2695 39028
rect 0 35187 125 39011
rect 2669 35187 2695 39011
rect 0 35186 2695 35187
rect 12301 39190 12306 39254
rect 12370 39190 12386 39254
rect 12450 39190 12466 39254
rect 12530 39190 12546 39254
rect 12610 39190 12626 39254
rect 12690 39190 12706 39254
rect 12770 39190 12786 39254
rect 12850 39190 12866 39254
rect 12930 39190 12946 39254
rect 13010 39190 13026 39254
rect 13090 39190 13106 39254
rect 13170 39190 13186 39254
rect 13250 39190 13266 39254
rect 13330 39190 13346 39254
rect 13410 39190 13426 39254
rect 13490 39190 13506 39254
rect 13570 39190 13586 39254
rect 13650 39190 13666 39254
rect 13730 39190 13746 39254
rect 13810 39190 13826 39254
rect 13890 39190 13906 39254
rect 13970 39190 13986 39254
rect 14050 39190 14066 39254
rect 14130 39190 14146 39254
rect 14210 39190 14226 39254
rect 14290 39190 14306 39254
rect 14370 39190 14386 39254
rect 14450 39190 14466 39254
rect 14530 39190 14546 39254
rect 14610 39190 14626 39254
rect 14690 39190 14706 39254
rect 14770 39190 14786 39254
rect 14850 39190 15000 39254
rect 12301 39173 15000 39190
rect 12301 39109 12306 39173
rect 12370 39109 12386 39173
rect 12450 39109 12466 39173
rect 12530 39109 12546 39173
rect 12610 39109 12626 39173
rect 12690 39109 12706 39173
rect 12770 39109 12786 39173
rect 12850 39109 12866 39173
rect 12930 39109 12946 39173
rect 13010 39109 13026 39173
rect 13090 39109 13106 39173
rect 13170 39109 13186 39173
rect 13250 39109 13266 39173
rect 13330 39109 13346 39173
rect 13410 39109 13426 39173
rect 13490 39109 13506 39173
rect 13570 39109 13586 39173
rect 13650 39109 13666 39173
rect 13730 39109 13746 39173
rect 13810 39109 13826 39173
rect 13890 39109 13906 39173
rect 13970 39109 13986 39173
rect 14050 39109 14066 39173
rect 14130 39109 14146 39173
rect 14210 39109 14226 39173
rect 14290 39109 14306 39173
rect 14370 39109 14386 39173
rect 14450 39109 14466 39173
rect 14530 39109 14546 39173
rect 14610 39109 14626 39173
rect 14690 39109 14706 39173
rect 14770 39109 14786 39173
rect 14850 39109 15000 39173
rect 12301 39092 15000 39109
rect 12301 39028 12306 39092
rect 12370 39028 12386 39092
rect 12450 39028 12466 39092
rect 12530 39028 12546 39092
rect 12610 39028 12626 39092
rect 12690 39028 12706 39092
rect 12770 39028 12786 39092
rect 12850 39028 12866 39092
rect 12930 39028 12946 39092
rect 13010 39028 13026 39092
rect 13090 39028 13106 39092
rect 13170 39028 13186 39092
rect 13250 39028 13266 39092
rect 13330 39028 13346 39092
rect 13410 39028 13426 39092
rect 13490 39028 13506 39092
rect 13570 39028 13586 39092
rect 13650 39028 13666 39092
rect 13730 39028 13746 39092
rect 13810 39028 13826 39092
rect 13890 39028 13906 39092
rect 13970 39028 13986 39092
rect 14050 39028 14066 39092
rect 14130 39028 14146 39092
rect 14210 39028 14226 39092
rect 14290 39028 14306 39092
rect 14370 39028 14386 39092
rect 14450 39028 14466 39092
rect 14530 39028 14546 39092
rect 14610 39028 14626 39092
rect 14690 39028 14706 39092
rect 14770 39028 14786 39092
rect 14850 39028 15000 39092
rect 12301 39011 15000 39028
rect 12301 35187 12306 39011
rect 14850 35187 15000 39011
rect 12301 35186 15000 35187
rect 0 35157 254 35186
rect 14746 35157 15000 35186
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 12534 4874 12537
rect 0 12470 105 12534
rect 169 12470 187 12534
rect 251 12470 269 12534
rect 333 12470 351 12534
rect 415 12470 433 12534
rect 497 12470 515 12534
rect 579 12470 597 12534
rect 661 12470 678 12534
rect 742 12470 759 12534
rect 823 12470 840 12534
rect 904 12470 921 12534
rect 985 12470 1002 12534
rect 1066 12470 1083 12534
rect 1147 12470 1164 12534
rect 1228 12470 1245 12534
rect 1309 12470 1326 12534
rect 1390 12470 1407 12534
rect 1471 12470 1488 12534
rect 1552 12470 1569 12534
rect 1633 12470 1650 12534
rect 1714 12470 1731 12534
rect 1795 12470 1812 12534
rect 1876 12470 1893 12534
rect 1957 12470 1974 12534
rect 2038 12470 2055 12534
rect 2119 12470 2136 12534
rect 2200 12470 2217 12534
rect 2281 12470 2298 12534
rect 2362 12470 2379 12534
rect 2443 12470 2460 12534
rect 2524 12470 2541 12534
rect 2605 12470 2622 12534
rect 2686 12470 2703 12534
rect 2767 12470 2784 12534
rect 2848 12470 2865 12534
rect 2929 12470 2946 12534
rect 3010 12470 3027 12534
rect 3091 12470 3108 12534
rect 3172 12470 3189 12534
rect 3253 12470 3270 12534
rect 3334 12470 3351 12534
rect 3415 12470 3432 12534
rect 3496 12470 3513 12534
rect 3577 12470 3594 12534
rect 3658 12470 3675 12534
rect 3739 12470 3756 12534
rect 3820 12470 3837 12534
rect 3901 12470 3918 12534
rect 3982 12470 3999 12534
rect 4063 12470 4080 12534
rect 4144 12470 4161 12534
rect 4225 12470 4242 12534
rect 4306 12470 4323 12534
rect 4387 12470 4404 12534
rect 4468 12470 4485 12534
rect 4549 12470 4566 12534
rect 4630 12470 4647 12534
rect 4711 12470 4728 12534
rect 4792 12470 4809 12534
rect 4873 12470 4874 12534
rect 0 12452 4874 12470
rect 0 12388 105 12452
rect 169 12388 187 12452
rect 251 12388 269 12452
rect 333 12388 351 12452
rect 415 12388 433 12452
rect 497 12388 515 12452
rect 579 12388 597 12452
rect 661 12388 678 12452
rect 742 12388 759 12452
rect 823 12388 840 12452
rect 904 12388 921 12452
rect 985 12388 1002 12452
rect 1066 12388 1083 12452
rect 1147 12388 1164 12452
rect 1228 12388 1245 12452
rect 1309 12388 1326 12452
rect 1390 12388 1407 12452
rect 1471 12388 1488 12452
rect 1552 12388 1569 12452
rect 1633 12388 1650 12452
rect 1714 12388 1731 12452
rect 1795 12388 1812 12452
rect 1876 12388 1893 12452
rect 1957 12388 1974 12452
rect 2038 12388 2055 12452
rect 2119 12388 2136 12452
rect 2200 12388 2217 12452
rect 2281 12388 2298 12452
rect 2362 12388 2379 12452
rect 2443 12388 2460 12452
rect 2524 12388 2541 12452
rect 2605 12388 2622 12452
rect 2686 12388 2703 12452
rect 2767 12388 2784 12452
rect 2848 12388 2865 12452
rect 2929 12388 2946 12452
rect 3010 12388 3027 12452
rect 3091 12388 3108 12452
rect 3172 12388 3189 12452
rect 3253 12388 3270 12452
rect 3334 12388 3351 12452
rect 3415 12388 3432 12452
rect 3496 12388 3513 12452
rect 3577 12388 3594 12452
rect 3658 12388 3675 12452
rect 3739 12388 3756 12452
rect 3820 12388 3837 12452
rect 3901 12388 3918 12452
rect 3982 12388 3999 12452
rect 4063 12388 4080 12452
rect 4144 12388 4161 12452
rect 4225 12388 4242 12452
rect 4306 12388 4323 12452
rect 4387 12388 4404 12452
rect 4468 12388 4485 12452
rect 4549 12388 4566 12452
rect 4630 12388 4647 12452
rect 4711 12388 4728 12452
rect 4792 12388 4809 12452
rect 4873 12388 4874 12452
rect 0 12370 4874 12388
rect 0 12306 105 12370
rect 169 12306 187 12370
rect 251 12306 269 12370
rect 333 12306 351 12370
rect 415 12306 433 12370
rect 497 12306 515 12370
rect 579 12306 597 12370
rect 661 12306 678 12370
rect 742 12306 759 12370
rect 823 12306 840 12370
rect 904 12306 921 12370
rect 985 12306 1002 12370
rect 1066 12306 1083 12370
rect 1147 12306 1164 12370
rect 1228 12306 1245 12370
rect 1309 12306 1326 12370
rect 1390 12306 1407 12370
rect 1471 12306 1488 12370
rect 1552 12306 1569 12370
rect 1633 12306 1650 12370
rect 1714 12306 1731 12370
rect 1795 12306 1812 12370
rect 1876 12306 1893 12370
rect 1957 12306 1974 12370
rect 2038 12306 2055 12370
rect 2119 12306 2136 12370
rect 2200 12306 2217 12370
rect 2281 12306 2298 12370
rect 2362 12306 2379 12370
rect 2443 12306 2460 12370
rect 2524 12306 2541 12370
rect 2605 12306 2622 12370
rect 2686 12306 2703 12370
rect 2767 12306 2784 12370
rect 2848 12306 2865 12370
rect 2929 12306 2946 12370
rect 3010 12306 3027 12370
rect 3091 12306 3108 12370
rect 3172 12306 3189 12370
rect 3253 12306 3270 12370
rect 3334 12306 3351 12370
rect 3415 12306 3432 12370
rect 3496 12306 3513 12370
rect 3577 12306 3594 12370
rect 3658 12306 3675 12370
rect 3739 12306 3756 12370
rect 3820 12306 3837 12370
rect 3901 12306 3918 12370
rect 3982 12306 3999 12370
rect 4063 12306 4080 12370
rect 4144 12306 4161 12370
rect 4225 12306 4242 12370
rect 4306 12306 4323 12370
rect 4387 12306 4404 12370
rect 4468 12306 4485 12370
rect 4549 12306 4566 12370
rect 4630 12306 4647 12370
rect 4711 12306 4728 12370
rect 4792 12306 4809 12370
rect 4873 12306 4874 12370
rect 0 12288 4874 12306
rect 0 12224 105 12288
rect 169 12224 187 12288
rect 251 12224 269 12288
rect 333 12224 351 12288
rect 415 12224 433 12288
rect 497 12224 515 12288
rect 579 12224 597 12288
rect 661 12224 678 12288
rect 742 12224 759 12288
rect 823 12224 840 12288
rect 904 12224 921 12288
rect 985 12224 1002 12288
rect 1066 12224 1083 12288
rect 1147 12224 1164 12288
rect 1228 12224 1245 12288
rect 1309 12224 1326 12288
rect 1390 12224 1407 12288
rect 1471 12224 1488 12288
rect 1552 12224 1569 12288
rect 1633 12224 1650 12288
rect 1714 12224 1731 12288
rect 1795 12224 1812 12288
rect 1876 12224 1893 12288
rect 1957 12224 1974 12288
rect 2038 12224 2055 12288
rect 2119 12224 2136 12288
rect 2200 12224 2217 12288
rect 2281 12224 2298 12288
rect 2362 12224 2379 12288
rect 2443 12224 2460 12288
rect 2524 12224 2541 12288
rect 2605 12224 2622 12288
rect 2686 12224 2703 12288
rect 2767 12224 2784 12288
rect 2848 12224 2865 12288
rect 2929 12224 2946 12288
rect 3010 12224 3027 12288
rect 3091 12224 3108 12288
rect 3172 12224 3189 12288
rect 3253 12224 3270 12288
rect 3334 12224 3351 12288
rect 3415 12224 3432 12288
rect 3496 12224 3513 12288
rect 3577 12224 3594 12288
rect 3658 12224 3675 12288
rect 3739 12224 3756 12288
rect 3820 12224 3837 12288
rect 3901 12224 3918 12288
rect 3982 12224 3999 12288
rect 4063 12224 4080 12288
rect 4144 12224 4161 12288
rect 4225 12224 4242 12288
rect 4306 12224 4323 12288
rect 4387 12224 4404 12288
rect 4468 12224 4485 12288
rect 4549 12224 4566 12288
rect 4630 12224 4647 12288
rect 4711 12224 4728 12288
rect 4792 12224 4809 12288
rect 4873 12224 4874 12288
rect 0 12206 4874 12224
rect 0 12142 105 12206
rect 169 12142 187 12206
rect 251 12142 269 12206
rect 333 12142 351 12206
rect 415 12142 433 12206
rect 497 12142 515 12206
rect 579 12142 597 12206
rect 661 12142 678 12206
rect 742 12142 759 12206
rect 823 12142 840 12206
rect 904 12142 921 12206
rect 985 12142 1002 12206
rect 1066 12142 1083 12206
rect 1147 12142 1164 12206
rect 1228 12142 1245 12206
rect 1309 12142 1326 12206
rect 1390 12142 1407 12206
rect 1471 12142 1488 12206
rect 1552 12142 1569 12206
rect 1633 12142 1650 12206
rect 1714 12142 1731 12206
rect 1795 12142 1812 12206
rect 1876 12142 1893 12206
rect 1957 12142 1974 12206
rect 2038 12142 2055 12206
rect 2119 12142 2136 12206
rect 2200 12142 2217 12206
rect 2281 12142 2298 12206
rect 2362 12142 2379 12206
rect 2443 12142 2460 12206
rect 2524 12142 2541 12206
rect 2605 12142 2622 12206
rect 2686 12142 2703 12206
rect 2767 12142 2784 12206
rect 2848 12142 2865 12206
rect 2929 12142 2946 12206
rect 3010 12142 3027 12206
rect 3091 12142 3108 12206
rect 3172 12142 3189 12206
rect 3253 12142 3270 12206
rect 3334 12142 3351 12206
rect 3415 12142 3432 12206
rect 3496 12142 3513 12206
rect 3577 12142 3594 12206
rect 3658 12142 3675 12206
rect 3739 12142 3756 12206
rect 3820 12142 3837 12206
rect 3901 12142 3918 12206
rect 3982 12142 3999 12206
rect 4063 12142 4080 12206
rect 4144 12142 4161 12206
rect 4225 12142 4242 12206
rect 4306 12142 4323 12206
rect 4387 12142 4404 12206
rect 4468 12142 4485 12206
rect 4549 12142 4566 12206
rect 4630 12142 4647 12206
rect 4711 12142 4728 12206
rect 4792 12142 4809 12206
rect 4873 12142 4874 12206
rect 0 12124 4874 12142
rect 0 12060 105 12124
rect 169 12060 187 12124
rect 251 12060 269 12124
rect 333 12060 351 12124
rect 415 12060 433 12124
rect 497 12060 515 12124
rect 579 12060 597 12124
rect 661 12060 678 12124
rect 742 12060 759 12124
rect 823 12060 840 12124
rect 904 12060 921 12124
rect 985 12060 1002 12124
rect 1066 12060 1083 12124
rect 1147 12060 1164 12124
rect 1228 12060 1245 12124
rect 1309 12060 1326 12124
rect 1390 12060 1407 12124
rect 1471 12060 1488 12124
rect 1552 12060 1569 12124
rect 1633 12060 1650 12124
rect 1714 12060 1731 12124
rect 1795 12060 1812 12124
rect 1876 12060 1893 12124
rect 1957 12060 1974 12124
rect 2038 12060 2055 12124
rect 2119 12060 2136 12124
rect 2200 12060 2217 12124
rect 2281 12060 2298 12124
rect 2362 12060 2379 12124
rect 2443 12060 2460 12124
rect 2524 12060 2541 12124
rect 2605 12060 2622 12124
rect 2686 12060 2703 12124
rect 2767 12060 2784 12124
rect 2848 12060 2865 12124
rect 2929 12060 2946 12124
rect 3010 12060 3027 12124
rect 3091 12060 3108 12124
rect 3172 12060 3189 12124
rect 3253 12060 3270 12124
rect 3334 12060 3351 12124
rect 3415 12060 3432 12124
rect 3496 12060 3513 12124
rect 3577 12060 3594 12124
rect 3658 12060 3675 12124
rect 3739 12060 3756 12124
rect 3820 12060 3837 12124
rect 3901 12060 3918 12124
rect 3982 12060 3999 12124
rect 4063 12060 4080 12124
rect 4144 12060 4161 12124
rect 4225 12060 4242 12124
rect 4306 12060 4323 12124
rect 4387 12060 4404 12124
rect 4468 12060 4485 12124
rect 4549 12060 4566 12124
rect 4630 12060 4647 12124
rect 4711 12060 4728 12124
rect 4792 12060 4809 12124
rect 4873 12060 4874 12124
rect 0 12042 4874 12060
rect 0 11978 105 12042
rect 169 11978 187 12042
rect 251 11978 269 12042
rect 333 11978 351 12042
rect 415 11978 433 12042
rect 497 11978 515 12042
rect 579 11978 597 12042
rect 661 11978 678 12042
rect 742 11978 759 12042
rect 823 11978 840 12042
rect 904 11978 921 12042
rect 985 11978 1002 12042
rect 1066 11978 1083 12042
rect 1147 11978 1164 12042
rect 1228 11978 1245 12042
rect 1309 11978 1326 12042
rect 1390 11978 1407 12042
rect 1471 11978 1488 12042
rect 1552 11978 1569 12042
rect 1633 11978 1650 12042
rect 1714 11978 1731 12042
rect 1795 11978 1812 12042
rect 1876 11978 1893 12042
rect 1957 11978 1974 12042
rect 2038 11978 2055 12042
rect 2119 11978 2136 12042
rect 2200 11978 2217 12042
rect 2281 11978 2298 12042
rect 2362 11978 2379 12042
rect 2443 11978 2460 12042
rect 2524 11978 2541 12042
rect 2605 11978 2622 12042
rect 2686 11978 2703 12042
rect 2767 11978 2784 12042
rect 2848 11978 2865 12042
rect 2929 11978 2946 12042
rect 3010 11978 3027 12042
rect 3091 11978 3108 12042
rect 3172 11978 3189 12042
rect 3253 11978 3270 12042
rect 3334 11978 3351 12042
rect 3415 11978 3432 12042
rect 3496 11978 3513 12042
rect 3577 11978 3594 12042
rect 3658 11978 3675 12042
rect 3739 11978 3756 12042
rect 3820 11978 3837 12042
rect 3901 11978 3918 12042
rect 3982 11978 3999 12042
rect 4063 11978 4080 12042
rect 4144 11978 4161 12042
rect 4225 11978 4242 12042
rect 4306 11978 4323 12042
rect 4387 11978 4404 12042
rect 4468 11978 4485 12042
rect 4549 11978 4566 12042
rect 4630 11978 4647 12042
rect 4711 11978 4728 12042
rect 4792 11978 4809 12042
rect 4873 11978 4874 12042
rect 0 11960 4874 11978
rect 0 11896 105 11960
rect 169 11896 187 11960
rect 251 11896 269 11960
rect 333 11896 351 11960
rect 415 11896 433 11960
rect 497 11896 515 11960
rect 579 11896 597 11960
rect 661 11896 678 11960
rect 742 11896 759 11960
rect 823 11896 840 11960
rect 904 11896 921 11960
rect 985 11896 1002 11960
rect 1066 11896 1083 11960
rect 1147 11896 1164 11960
rect 1228 11896 1245 11960
rect 1309 11896 1326 11960
rect 1390 11896 1407 11960
rect 1471 11896 1488 11960
rect 1552 11896 1569 11960
rect 1633 11896 1650 11960
rect 1714 11896 1731 11960
rect 1795 11896 1812 11960
rect 1876 11896 1893 11960
rect 1957 11896 1974 11960
rect 2038 11896 2055 11960
rect 2119 11896 2136 11960
rect 2200 11896 2217 11960
rect 2281 11896 2298 11960
rect 2362 11896 2379 11960
rect 2443 11896 2460 11960
rect 2524 11896 2541 11960
rect 2605 11896 2622 11960
rect 2686 11896 2703 11960
rect 2767 11896 2784 11960
rect 2848 11896 2865 11960
rect 2929 11896 2946 11960
rect 3010 11896 3027 11960
rect 3091 11896 3108 11960
rect 3172 11896 3189 11960
rect 3253 11896 3270 11960
rect 3334 11896 3351 11960
rect 3415 11896 3432 11960
rect 3496 11896 3513 11960
rect 3577 11896 3594 11960
rect 3658 11896 3675 11960
rect 3739 11896 3756 11960
rect 3820 11896 3837 11960
rect 3901 11896 3918 11960
rect 3982 11896 3999 11960
rect 4063 11896 4080 11960
rect 4144 11896 4161 11960
rect 4225 11896 4242 11960
rect 4306 11896 4323 11960
rect 4387 11896 4404 11960
rect 4468 11896 4485 11960
rect 4549 11896 4566 11960
rect 4630 11896 4647 11960
rect 4711 11896 4728 11960
rect 4792 11896 4809 11960
rect 4873 11896 4874 11960
rect 0 11878 4874 11896
rect 0 11814 105 11878
rect 169 11814 187 11878
rect 251 11814 269 11878
rect 333 11814 351 11878
rect 415 11814 433 11878
rect 497 11814 515 11878
rect 579 11814 597 11878
rect 661 11814 678 11878
rect 742 11814 759 11878
rect 823 11814 840 11878
rect 904 11814 921 11878
rect 985 11814 1002 11878
rect 1066 11814 1083 11878
rect 1147 11814 1164 11878
rect 1228 11814 1245 11878
rect 1309 11814 1326 11878
rect 1390 11814 1407 11878
rect 1471 11814 1488 11878
rect 1552 11814 1569 11878
rect 1633 11814 1650 11878
rect 1714 11814 1731 11878
rect 1795 11814 1812 11878
rect 1876 11814 1893 11878
rect 1957 11814 1974 11878
rect 2038 11814 2055 11878
rect 2119 11814 2136 11878
rect 2200 11814 2217 11878
rect 2281 11814 2298 11878
rect 2362 11814 2379 11878
rect 2443 11814 2460 11878
rect 2524 11814 2541 11878
rect 2605 11814 2622 11878
rect 2686 11814 2703 11878
rect 2767 11814 2784 11878
rect 2848 11814 2865 11878
rect 2929 11814 2946 11878
rect 3010 11814 3027 11878
rect 3091 11814 3108 11878
rect 3172 11814 3189 11878
rect 3253 11814 3270 11878
rect 3334 11814 3351 11878
rect 3415 11814 3432 11878
rect 3496 11814 3513 11878
rect 3577 11814 3594 11878
rect 3658 11814 3675 11878
rect 3739 11814 3756 11878
rect 3820 11814 3837 11878
rect 3901 11814 3918 11878
rect 3982 11814 3999 11878
rect 4063 11814 4080 11878
rect 4144 11814 4161 11878
rect 4225 11814 4242 11878
rect 4306 11814 4323 11878
rect 4387 11814 4404 11878
rect 4468 11814 4485 11878
rect 4549 11814 4566 11878
rect 4630 11814 4647 11878
rect 4711 11814 4728 11878
rect 4792 11814 4809 11878
rect 4873 11814 4874 11878
rect 0 11796 4874 11814
rect 0 11732 105 11796
rect 169 11732 187 11796
rect 251 11732 269 11796
rect 333 11732 351 11796
rect 415 11732 433 11796
rect 497 11732 515 11796
rect 579 11732 597 11796
rect 661 11732 678 11796
rect 742 11732 759 11796
rect 823 11732 840 11796
rect 904 11732 921 11796
rect 985 11732 1002 11796
rect 1066 11732 1083 11796
rect 1147 11732 1164 11796
rect 1228 11732 1245 11796
rect 1309 11732 1326 11796
rect 1390 11732 1407 11796
rect 1471 11732 1488 11796
rect 1552 11732 1569 11796
rect 1633 11732 1650 11796
rect 1714 11732 1731 11796
rect 1795 11732 1812 11796
rect 1876 11732 1893 11796
rect 1957 11732 1974 11796
rect 2038 11732 2055 11796
rect 2119 11732 2136 11796
rect 2200 11732 2217 11796
rect 2281 11732 2298 11796
rect 2362 11732 2379 11796
rect 2443 11732 2460 11796
rect 2524 11732 2541 11796
rect 2605 11732 2622 11796
rect 2686 11732 2703 11796
rect 2767 11732 2784 11796
rect 2848 11732 2865 11796
rect 2929 11732 2946 11796
rect 3010 11732 3027 11796
rect 3091 11732 3108 11796
rect 3172 11732 3189 11796
rect 3253 11732 3270 11796
rect 3334 11732 3351 11796
rect 3415 11732 3432 11796
rect 3496 11732 3513 11796
rect 3577 11732 3594 11796
rect 3658 11732 3675 11796
rect 3739 11732 3756 11796
rect 3820 11732 3837 11796
rect 3901 11732 3918 11796
rect 3982 11732 3999 11796
rect 4063 11732 4080 11796
rect 4144 11732 4161 11796
rect 4225 11732 4242 11796
rect 4306 11732 4323 11796
rect 4387 11732 4404 11796
rect 4468 11732 4485 11796
rect 4549 11732 4566 11796
rect 4630 11732 4647 11796
rect 4711 11732 4728 11796
rect 4792 11732 4809 11796
rect 4873 11732 4874 11796
rect 0 11714 4874 11732
rect 0 11650 105 11714
rect 169 11650 187 11714
rect 251 11650 269 11714
rect 333 11650 351 11714
rect 415 11650 433 11714
rect 497 11650 515 11714
rect 579 11650 597 11714
rect 661 11650 678 11714
rect 742 11650 759 11714
rect 823 11650 840 11714
rect 904 11650 921 11714
rect 985 11650 1002 11714
rect 1066 11650 1083 11714
rect 1147 11650 1164 11714
rect 1228 11650 1245 11714
rect 1309 11650 1326 11714
rect 1390 11650 1407 11714
rect 1471 11650 1488 11714
rect 1552 11650 1569 11714
rect 1633 11650 1650 11714
rect 1714 11650 1731 11714
rect 1795 11650 1812 11714
rect 1876 11650 1893 11714
rect 1957 11650 1974 11714
rect 2038 11650 2055 11714
rect 2119 11650 2136 11714
rect 2200 11650 2217 11714
rect 2281 11650 2298 11714
rect 2362 11650 2379 11714
rect 2443 11650 2460 11714
rect 2524 11650 2541 11714
rect 2605 11650 2622 11714
rect 2686 11650 2703 11714
rect 2767 11650 2784 11714
rect 2848 11650 2865 11714
rect 2929 11650 2946 11714
rect 3010 11650 3027 11714
rect 3091 11650 3108 11714
rect 3172 11650 3189 11714
rect 3253 11650 3270 11714
rect 3334 11650 3351 11714
rect 3415 11650 3432 11714
rect 3496 11650 3513 11714
rect 3577 11650 3594 11714
rect 3658 11650 3675 11714
rect 3739 11650 3756 11714
rect 3820 11650 3837 11714
rect 3901 11650 3918 11714
rect 3982 11650 3999 11714
rect 4063 11650 4080 11714
rect 4144 11650 4161 11714
rect 4225 11650 4242 11714
rect 4306 11650 4323 11714
rect 4387 11650 4404 11714
rect 4468 11650 4485 11714
rect 4549 11650 4566 11714
rect 4630 11650 4647 11714
rect 4711 11650 4728 11714
rect 4792 11650 4809 11714
rect 4873 11650 4874 11714
rect 0 11647 4874 11650
rect 10083 12534 15000 12537
rect 10083 12470 10084 12534
rect 10148 12470 10166 12534
rect 10230 12470 10248 12534
rect 10312 12470 10330 12534
rect 10394 12470 10412 12534
rect 10476 12470 10494 12534
rect 10558 12470 10576 12534
rect 10640 12470 10657 12534
rect 10721 12470 10738 12534
rect 10802 12470 10819 12534
rect 10883 12470 10900 12534
rect 10964 12470 10981 12534
rect 11045 12470 11062 12534
rect 11126 12470 11143 12534
rect 11207 12470 11224 12534
rect 11288 12470 11305 12534
rect 11369 12470 11386 12534
rect 11450 12470 11467 12534
rect 11531 12470 11548 12534
rect 11612 12470 11629 12534
rect 11693 12470 11710 12534
rect 11774 12470 11791 12534
rect 11855 12470 11872 12534
rect 11936 12470 11953 12534
rect 12017 12470 12034 12534
rect 12098 12470 12115 12534
rect 12179 12470 12196 12534
rect 12260 12470 12277 12534
rect 12341 12470 12358 12534
rect 12422 12470 12439 12534
rect 12503 12470 12520 12534
rect 12584 12470 12601 12534
rect 12665 12470 12682 12534
rect 12746 12470 12763 12534
rect 12827 12470 12844 12534
rect 12908 12470 12925 12534
rect 12989 12470 13006 12534
rect 13070 12470 13087 12534
rect 13151 12470 13168 12534
rect 13232 12470 13249 12534
rect 13313 12470 13330 12534
rect 13394 12470 13411 12534
rect 13475 12470 13492 12534
rect 13556 12470 13573 12534
rect 13637 12470 13654 12534
rect 13718 12470 13735 12534
rect 13799 12470 13816 12534
rect 13880 12470 13897 12534
rect 13961 12470 13978 12534
rect 14042 12470 14059 12534
rect 14123 12470 14140 12534
rect 14204 12470 14221 12534
rect 14285 12470 14302 12534
rect 14366 12470 14383 12534
rect 14447 12470 14464 12534
rect 14528 12470 14545 12534
rect 14609 12470 14626 12534
rect 14690 12470 14707 12534
rect 14771 12470 14788 12534
rect 14852 12470 15000 12534
rect 10083 12452 15000 12470
rect 10083 12388 10084 12452
rect 10148 12388 10166 12452
rect 10230 12388 10248 12452
rect 10312 12388 10330 12452
rect 10394 12388 10412 12452
rect 10476 12388 10494 12452
rect 10558 12388 10576 12452
rect 10640 12388 10657 12452
rect 10721 12388 10738 12452
rect 10802 12388 10819 12452
rect 10883 12388 10900 12452
rect 10964 12388 10981 12452
rect 11045 12388 11062 12452
rect 11126 12388 11143 12452
rect 11207 12388 11224 12452
rect 11288 12388 11305 12452
rect 11369 12388 11386 12452
rect 11450 12388 11467 12452
rect 11531 12388 11548 12452
rect 11612 12388 11629 12452
rect 11693 12388 11710 12452
rect 11774 12388 11791 12452
rect 11855 12388 11872 12452
rect 11936 12388 11953 12452
rect 12017 12388 12034 12452
rect 12098 12388 12115 12452
rect 12179 12388 12196 12452
rect 12260 12388 12277 12452
rect 12341 12388 12358 12452
rect 12422 12388 12439 12452
rect 12503 12388 12520 12452
rect 12584 12388 12601 12452
rect 12665 12388 12682 12452
rect 12746 12388 12763 12452
rect 12827 12388 12844 12452
rect 12908 12388 12925 12452
rect 12989 12388 13006 12452
rect 13070 12388 13087 12452
rect 13151 12388 13168 12452
rect 13232 12388 13249 12452
rect 13313 12388 13330 12452
rect 13394 12388 13411 12452
rect 13475 12388 13492 12452
rect 13556 12388 13573 12452
rect 13637 12388 13654 12452
rect 13718 12388 13735 12452
rect 13799 12388 13816 12452
rect 13880 12388 13897 12452
rect 13961 12388 13978 12452
rect 14042 12388 14059 12452
rect 14123 12388 14140 12452
rect 14204 12388 14221 12452
rect 14285 12388 14302 12452
rect 14366 12388 14383 12452
rect 14447 12388 14464 12452
rect 14528 12388 14545 12452
rect 14609 12388 14626 12452
rect 14690 12388 14707 12452
rect 14771 12388 14788 12452
rect 14852 12388 15000 12452
rect 10083 12370 15000 12388
rect 10083 12306 10084 12370
rect 10148 12306 10166 12370
rect 10230 12306 10248 12370
rect 10312 12306 10330 12370
rect 10394 12306 10412 12370
rect 10476 12306 10494 12370
rect 10558 12306 10576 12370
rect 10640 12306 10657 12370
rect 10721 12306 10738 12370
rect 10802 12306 10819 12370
rect 10883 12306 10900 12370
rect 10964 12306 10981 12370
rect 11045 12306 11062 12370
rect 11126 12306 11143 12370
rect 11207 12306 11224 12370
rect 11288 12306 11305 12370
rect 11369 12306 11386 12370
rect 11450 12306 11467 12370
rect 11531 12306 11548 12370
rect 11612 12306 11629 12370
rect 11693 12306 11710 12370
rect 11774 12306 11791 12370
rect 11855 12306 11872 12370
rect 11936 12306 11953 12370
rect 12017 12306 12034 12370
rect 12098 12306 12115 12370
rect 12179 12306 12196 12370
rect 12260 12306 12277 12370
rect 12341 12306 12358 12370
rect 12422 12306 12439 12370
rect 12503 12306 12520 12370
rect 12584 12306 12601 12370
rect 12665 12306 12682 12370
rect 12746 12306 12763 12370
rect 12827 12306 12844 12370
rect 12908 12306 12925 12370
rect 12989 12306 13006 12370
rect 13070 12306 13087 12370
rect 13151 12306 13168 12370
rect 13232 12306 13249 12370
rect 13313 12306 13330 12370
rect 13394 12306 13411 12370
rect 13475 12306 13492 12370
rect 13556 12306 13573 12370
rect 13637 12306 13654 12370
rect 13718 12306 13735 12370
rect 13799 12306 13816 12370
rect 13880 12306 13897 12370
rect 13961 12306 13978 12370
rect 14042 12306 14059 12370
rect 14123 12306 14140 12370
rect 14204 12306 14221 12370
rect 14285 12306 14302 12370
rect 14366 12306 14383 12370
rect 14447 12306 14464 12370
rect 14528 12306 14545 12370
rect 14609 12306 14626 12370
rect 14690 12306 14707 12370
rect 14771 12306 14788 12370
rect 14852 12306 15000 12370
rect 10083 12288 15000 12306
rect 10083 12224 10084 12288
rect 10148 12224 10166 12288
rect 10230 12224 10248 12288
rect 10312 12224 10330 12288
rect 10394 12224 10412 12288
rect 10476 12224 10494 12288
rect 10558 12224 10576 12288
rect 10640 12224 10657 12288
rect 10721 12224 10738 12288
rect 10802 12224 10819 12288
rect 10883 12224 10900 12288
rect 10964 12224 10981 12288
rect 11045 12224 11062 12288
rect 11126 12224 11143 12288
rect 11207 12224 11224 12288
rect 11288 12224 11305 12288
rect 11369 12224 11386 12288
rect 11450 12224 11467 12288
rect 11531 12224 11548 12288
rect 11612 12224 11629 12288
rect 11693 12224 11710 12288
rect 11774 12224 11791 12288
rect 11855 12224 11872 12288
rect 11936 12224 11953 12288
rect 12017 12224 12034 12288
rect 12098 12224 12115 12288
rect 12179 12224 12196 12288
rect 12260 12224 12277 12288
rect 12341 12224 12358 12288
rect 12422 12224 12439 12288
rect 12503 12224 12520 12288
rect 12584 12224 12601 12288
rect 12665 12224 12682 12288
rect 12746 12224 12763 12288
rect 12827 12224 12844 12288
rect 12908 12224 12925 12288
rect 12989 12224 13006 12288
rect 13070 12224 13087 12288
rect 13151 12224 13168 12288
rect 13232 12224 13249 12288
rect 13313 12224 13330 12288
rect 13394 12224 13411 12288
rect 13475 12224 13492 12288
rect 13556 12224 13573 12288
rect 13637 12224 13654 12288
rect 13718 12224 13735 12288
rect 13799 12224 13816 12288
rect 13880 12224 13897 12288
rect 13961 12224 13978 12288
rect 14042 12224 14059 12288
rect 14123 12224 14140 12288
rect 14204 12224 14221 12288
rect 14285 12224 14302 12288
rect 14366 12224 14383 12288
rect 14447 12224 14464 12288
rect 14528 12224 14545 12288
rect 14609 12224 14626 12288
rect 14690 12224 14707 12288
rect 14771 12224 14788 12288
rect 14852 12224 15000 12288
rect 10083 12206 15000 12224
rect 10083 12142 10084 12206
rect 10148 12142 10166 12206
rect 10230 12142 10248 12206
rect 10312 12142 10330 12206
rect 10394 12142 10412 12206
rect 10476 12142 10494 12206
rect 10558 12142 10576 12206
rect 10640 12142 10657 12206
rect 10721 12142 10738 12206
rect 10802 12142 10819 12206
rect 10883 12142 10900 12206
rect 10964 12142 10981 12206
rect 11045 12142 11062 12206
rect 11126 12142 11143 12206
rect 11207 12142 11224 12206
rect 11288 12142 11305 12206
rect 11369 12142 11386 12206
rect 11450 12142 11467 12206
rect 11531 12142 11548 12206
rect 11612 12142 11629 12206
rect 11693 12142 11710 12206
rect 11774 12142 11791 12206
rect 11855 12142 11872 12206
rect 11936 12142 11953 12206
rect 12017 12142 12034 12206
rect 12098 12142 12115 12206
rect 12179 12142 12196 12206
rect 12260 12142 12277 12206
rect 12341 12142 12358 12206
rect 12422 12142 12439 12206
rect 12503 12142 12520 12206
rect 12584 12142 12601 12206
rect 12665 12142 12682 12206
rect 12746 12142 12763 12206
rect 12827 12142 12844 12206
rect 12908 12142 12925 12206
rect 12989 12142 13006 12206
rect 13070 12142 13087 12206
rect 13151 12142 13168 12206
rect 13232 12142 13249 12206
rect 13313 12142 13330 12206
rect 13394 12142 13411 12206
rect 13475 12142 13492 12206
rect 13556 12142 13573 12206
rect 13637 12142 13654 12206
rect 13718 12142 13735 12206
rect 13799 12142 13816 12206
rect 13880 12142 13897 12206
rect 13961 12142 13978 12206
rect 14042 12142 14059 12206
rect 14123 12142 14140 12206
rect 14204 12142 14221 12206
rect 14285 12142 14302 12206
rect 14366 12142 14383 12206
rect 14447 12142 14464 12206
rect 14528 12142 14545 12206
rect 14609 12142 14626 12206
rect 14690 12142 14707 12206
rect 14771 12142 14788 12206
rect 14852 12142 15000 12206
rect 10083 12124 15000 12142
rect 10083 12060 10084 12124
rect 10148 12060 10166 12124
rect 10230 12060 10248 12124
rect 10312 12060 10330 12124
rect 10394 12060 10412 12124
rect 10476 12060 10494 12124
rect 10558 12060 10576 12124
rect 10640 12060 10657 12124
rect 10721 12060 10738 12124
rect 10802 12060 10819 12124
rect 10883 12060 10900 12124
rect 10964 12060 10981 12124
rect 11045 12060 11062 12124
rect 11126 12060 11143 12124
rect 11207 12060 11224 12124
rect 11288 12060 11305 12124
rect 11369 12060 11386 12124
rect 11450 12060 11467 12124
rect 11531 12060 11548 12124
rect 11612 12060 11629 12124
rect 11693 12060 11710 12124
rect 11774 12060 11791 12124
rect 11855 12060 11872 12124
rect 11936 12060 11953 12124
rect 12017 12060 12034 12124
rect 12098 12060 12115 12124
rect 12179 12060 12196 12124
rect 12260 12060 12277 12124
rect 12341 12060 12358 12124
rect 12422 12060 12439 12124
rect 12503 12060 12520 12124
rect 12584 12060 12601 12124
rect 12665 12060 12682 12124
rect 12746 12060 12763 12124
rect 12827 12060 12844 12124
rect 12908 12060 12925 12124
rect 12989 12060 13006 12124
rect 13070 12060 13087 12124
rect 13151 12060 13168 12124
rect 13232 12060 13249 12124
rect 13313 12060 13330 12124
rect 13394 12060 13411 12124
rect 13475 12060 13492 12124
rect 13556 12060 13573 12124
rect 13637 12060 13654 12124
rect 13718 12060 13735 12124
rect 13799 12060 13816 12124
rect 13880 12060 13897 12124
rect 13961 12060 13978 12124
rect 14042 12060 14059 12124
rect 14123 12060 14140 12124
rect 14204 12060 14221 12124
rect 14285 12060 14302 12124
rect 14366 12060 14383 12124
rect 14447 12060 14464 12124
rect 14528 12060 14545 12124
rect 14609 12060 14626 12124
rect 14690 12060 14707 12124
rect 14771 12060 14788 12124
rect 14852 12060 15000 12124
rect 10083 12042 15000 12060
rect 10083 11978 10084 12042
rect 10148 11978 10166 12042
rect 10230 11978 10248 12042
rect 10312 11978 10330 12042
rect 10394 11978 10412 12042
rect 10476 11978 10494 12042
rect 10558 11978 10576 12042
rect 10640 11978 10657 12042
rect 10721 11978 10738 12042
rect 10802 11978 10819 12042
rect 10883 11978 10900 12042
rect 10964 11978 10981 12042
rect 11045 11978 11062 12042
rect 11126 11978 11143 12042
rect 11207 11978 11224 12042
rect 11288 11978 11305 12042
rect 11369 11978 11386 12042
rect 11450 11978 11467 12042
rect 11531 11978 11548 12042
rect 11612 11978 11629 12042
rect 11693 11978 11710 12042
rect 11774 11978 11791 12042
rect 11855 11978 11872 12042
rect 11936 11978 11953 12042
rect 12017 11978 12034 12042
rect 12098 11978 12115 12042
rect 12179 11978 12196 12042
rect 12260 11978 12277 12042
rect 12341 11978 12358 12042
rect 12422 11978 12439 12042
rect 12503 11978 12520 12042
rect 12584 11978 12601 12042
rect 12665 11978 12682 12042
rect 12746 11978 12763 12042
rect 12827 11978 12844 12042
rect 12908 11978 12925 12042
rect 12989 11978 13006 12042
rect 13070 11978 13087 12042
rect 13151 11978 13168 12042
rect 13232 11978 13249 12042
rect 13313 11978 13330 12042
rect 13394 11978 13411 12042
rect 13475 11978 13492 12042
rect 13556 11978 13573 12042
rect 13637 11978 13654 12042
rect 13718 11978 13735 12042
rect 13799 11978 13816 12042
rect 13880 11978 13897 12042
rect 13961 11978 13978 12042
rect 14042 11978 14059 12042
rect 14123 11978 14140 12042
rect 14204 11978 14221 12042
rect 14285 11978 14302 12042
rect 14366 11978 14383 12042
rect 14447 11978 14464 12042
rect 14528 11978 14545 12042
rect 14609 11978 14626 12042
rect 14690 11978 14707 12042
rect 14771 11978 14788 12042
rect 14852 11978 15000 12042
rect 10083 11960 15000 11978
rect 10083 11896 10084 11960
rect 10148 11896 10166 11960
rect 10230 11896 10248 11960
rect 10312 11896 10330 11960
rect 10394 11896 10412 11960
rect 10476 11896 10494 11960
rect 10558 11896 10576 11960
rect 10640 11896 10657 11960
rect 10721 11896 10738 11960
rect 10802 11896 10819 11960
rect 10883 11896 10900 11960
rect 10964 11896 10981 11960
rect 11045 11896 11062 11960
rect 11126 11896 11143 11960
rect 11207 11896 11224 11960
rect 11288 11896 11305 11960
rect 11369 11896 11386 11960
rect 11450 11896 11467 11960
rect 11531 11896 11548 11960
rect 11612 11896 11629 11960
rect 11693 11896 11710 11960
rect 11774 11896 11791 11960
rect 11855 11896 11872 11960
rect 11936 11896 11953 11960
rect 12017 11896 12034 11960
rect 12098 11896 12115 11960
rect 12179 11896 12196 11960
rect 12260 11896 12277 11960
rect 12341 11896 12358 11960
rect 12422 11896 12439 11960
rect 12503 11896 12520 11960
rect 12584 11896 12601 11960
rect 12665 11896 12682 11960
rect 12746 11896 12763 11960
rect 12827 11896 12844 11960
rect 12908 11896 12925 11960
rect 12989 11896 13006 11960
rect 13070 11896 13087 11960
rect 13151 11896 13168 11960
rect 13232 11896 13249 11960
rect 13313 11896 13330 11960
rect 13394 11896 13411 11960
rect 13475 11896 13492 11960
rect 13556 11896 13573 11960
rect 13637 11896 13654 11960
rect 13718 11896 13735 11960
rect 13799 11896 13816 11960
rect 13880 11896 13897 11960
rect 13961 11896 13978 11960
rect 14042 11896 14059 11960
rect 14123 11896 14140 11960
rect 14204 11896 14221 11960
rect 14285 11896 14302 11960
rect 14366 11896 14383 11960
rect 14447 11896 14464 11960
rect 14528 11896 14545 11960
rect 14609 11896 14626 11960
rect 14690 11896 14707 11960
rect 14771 11896 14788 11960
rect 14852 11896 15000 11960
rect 10083 11878 15000 11896
rect 10083 11814 10084 11878
rect 10148 11814 10166 11878
rect 10230 11814 10248 11878
rect 10312 11814 10330 11878
rect 10394 11814 10412 11878
rect 10476 11814 10494 11878
rect 10558 11814 10576 11878
rect 10640 11814 10657 11878
rect 10721 11814 10738 11878
rect 10802 11814 10819 11878
rect 10883 11814 10900 11878
rect 10964 11814 10981 11878
rect 11045 11814 11062 11878
rect 11126 11814 11143 11878
rect 11207 11814 11224 11878
rect 11288 11814 11305 11878
rect 11369 11814 11386 11878
rect 11450 11814 11467 11878
rect 11531 11814 11548 11878
rect 11612 11814 11629 11878
rect 11693 11814 11710 11878
rect 11774 11814 11791 11878
rect 11855 11814 11872 11878
rect 11936 11814 11953 11878
rect 12017 11814 12034 11878
rect 12098 11814 12115 11878
rect 12179 11814 12196 11878
rect 12260 11814 12277 11878
rect 12341 11814 12358 11878
rect 12422 11814 12439 11878
rect 12503 11814 12520 11878
rect 12584 11814 12601 11878
rect 12665 11814 12682 11878
rect 12746 11814 12763 11878
rect 12827 11814 12844 11878
rect 12908 11814 12925 11878
rect 12989 11814 13006 11878
rect 13070 11814 13087 11878
rect 13151 11814 13168 11878
rect 13232 11814 13249 11878
rect 13313 11814 13330 11878
rect 13394 11814 13411 11878
rect 13475 11814 13492 11878
rect 13556 11814 13573 11878
rect 13637 11814 13654 11878
rect 13718 11814 13735 11878
rect 13799 11814 13816 11878
rect 13880 11814 13897 11878
rect 13961 11814 13978 11878
rect 14042 11814 14059 11878
rect 14123 11814 14140 11878
rect 14204 11814 14221 11878
rect 14285 11814 14302 11878
rect 14366 11814 14383 11878
rect 14447 11814 14464 11878
rect 14528 11814 14545 11878
rect 14609 11814 14626 11878
rect 14690 11814 14707 11878
rect 14771 11814 14788 11878
rect 14852 11814 15000 11878
rect 10083 11796 15000 11814
rect 10083 11732 10084 11796
rect 10148 11732 10166 11796
rect 10230 11732 10248 11796
rect 10312 11732 10330 11796
rect 10394 11732 10412 11796
rect 10476 11732 10494 11796
rect 10558 11732 10576 11796
rect 10640 11732 10657 11796
rect 10721 11732 10738 11796
rect 10802 11732 10819 11796
rect 10883 11732 10900 11796
rect 10964 11732 10981 11796
rect 11045 11732 11062 11796
rect 11126 11732 11143 11796
rect 11207 11732 11224 11796
rect 11288 11732 11305 11796
rect 11369 11732 11386 11796
rect 11450 11732 11467 11796
rect 11531 11732 11548 11796
rect 11612 11732 11629 11796
rect 11693 11732 11710 11796
rect 11774 11732 11791 11796
rect 11855 11732 11872 11796
rect 11936 11732 11953 11796
rect 12017 11732 12034 11796
rect 12098 11732 12115 11796
rect 12179 11732 12196 11796
rect 12260 11732 12277 11796
rect 12341 11732 12358 11796
rect 12422 11732 12439 11796
rect 12503 11732 12520 11796
rect 12584 11732 12601 11796
rect 12665 11732 12682 11796
rect 12746 11732 12763 11796
rect 12827 11732 12844 11796
rect 12908 11732 12925 11796
rect 12989 11732 13006 11796
rect 13070 11732 13087 11796
rect 13151 11732 13168 11796
rect 13232 11732 13249 11796
rect 13313 11732 13330 11796
rect 13394 11732 13411 11796
rect 13475 11732 13492 11796
rect 13556 11732 13573 11796
rect 13637 11732 13654 11796
rect 13718 11732 13735 11796
rect 13799 11732 13816 11796
rect 13880 11732 13897 11796
rect 13961 11732 13978 11796
rect 14042 11732 14059 11796
rect 14123 11732 14140 11796
rect 14204 11732 14221 11796
rect 14285 11732 14302 11796
rect 14366 11732 14383 11796
rect 14447 11732 14464 11796
rect 14528 11732 14545 11796
rect 14609 11732 14626 11796
rect 14690 11732 14707 11796
rect 14771 11732 14788 11796
rect 14852 11732 15000 11796
rect 10083 11714 15000 11732
rect 10083 11650 10084 11714
rect 10148 11650 10166 11714
rect 10230 11650 10248 11714
rect 10312 11650 10330 11714
rect 10394 11650 10412 11714
rect 10476 11650 10494 11714
rect 10558 11650 10576 11714
rect 10640 11650 10657 11714
rect 10721 11650 10738 11714
rect 10802 11650 10819 11714
rect 10883 11650 10900 11714
rect 10964 11650 10981 11714
rect 11045 11650 11062 11714
rect 11126 11650 11143 11714
rect 11207 11650 11224 11714
rect 11288 11650 11305 11714
rect 11369 11650 11386 11714
rect 11450 11650 11467 11714
rect 11531 11650 11548 11714
rect 11612 11650 11629 11714
rect 11693 11650 11710 11714
rect 11774 11650 11791 11714
rect 11855 11650 11872 11714
rect 11936 11650 11953 11714
rect 12017 11650 12034 11714
rect 12098 11650 12115 11714
rect 12179 11650 12196 11714
rect 12260 11650 12277 11714
rect 12341 11650 12358 11714
rect 12422 11650 12439 11714
rect 12503 11650 12520 11714
rect 12584 11650 12601 11714
rect 12665 11650 12682 11714
rect 12746 11650 12763 11714
rect 12827 11650 12844 11714
rect 12908 11650 12925 11714
rect 12989 11650 13006 11714
rect 13070 11650 13087 11714
rect 13151 11650 13168 11714
rect 13232 11650 13249 11714
rect 13313 11650 13330 11714
rect 13394 11650 13411 11714
rect 13475 11650 13492 11714
rect 13556 11650 13573 11714
rect 13637 11650 13654 11714
rect 13718 11650 13735 11714
rect 13799 11650 13816 11714
rect 13880 11650 13897 11714
rect 13961 11650 13978 11714
rect 14042 11650 14059 11714
rect 14123 11650 14140 11714
rect 14204 11650 14221 11714
rect 14285 11650 14302 11714
rect 14366 11650 14383 11714
rect 14447 11650 14464 11714
rect 14528 11650 14545 11714
rect 14609 11650 14626 11714
rect 14690 11650 14707 11714
rect 14771 11650 14788 11714
rect 14852 11650 15000 11714
rect 10083 11647 15000 11650
rect 0 11281 254 11347
rect 14746 11281 15000 11347
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9547 254 9613
rect 14746 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 6094 4874 6097
rect 0 6030 105 6094
rect 169 6030 187 6094
rect 251 6030 269 6094
rect 333 6030 351 6094
rect 415 6030 433 6094
rect 497 6030 515 6094
rect 579 6030 597 6094
rect 661 6030 678 6094
rect 742 6030 759 6094
rect 823 6030 840 6094
rect 904 6030 921 6094
rect 985 6030 1002 6094
rect 1066 6030 1083 6094
rect 1147 6030 1164 6094
rect 1228 6030 1245 6094
rect 1309 6030 1326 6094
rect 1390 6030 1407 6094
rect 1471 6030 1488 6094
rect 1552 6030 1569 6094
rect 1633 6030 1650 6094
rect 1714 6030 1731 6094
rect 1795 6030 1812 6094
rect 1876 6030 1893 6094
rect 1957 6030 1974 6094
rect 2038 6030 2055 6094
rect 2119 6030 2136 6094
rect 2200 6030 2217 6094
rect 2281 6030 2298 6094
rect 2362 6030 2379 6094
rect 2443 6030 2460 6094
rect 2524 6030 2541 6094
rect 2605 6030 2622 6094
rect 2686 6030 2703 6094
rect 2767 6030 2784 6094
rect 2848 6030 2865 6094
rect 2929 6030 2946 6094
rect 3010 6030 3027 6094
rect 3091 6030 3108 6094
rect 3172 6030 3189 6094
rect 3253 6030 3270 6094
rect 3334 6030 3351 6094
rect 3415 6030 3432 6094
rect 3496 6030 3513 6094
rect 3577 6030 3594 6094
rect 3658 6030 3675 6094
rect 3739 6030 3756 6094
rect 3820 6030 3837 6094
rect 3901 6030 3918 6094
rect 3982 6030 3999 6094
rect 4063 6030 4080 6094
rect 4144 6030 4161 6094
rect 4225 6030 4242 6094
rect 4306 6030 4323 6094
rect 4387 6030 4404 6094
rect 4468 6030 4485 6094
rect 4549 6030 4566 6094
rect 4630 6030 4647 6094
rect 4711 6030 4728 6094
rect 4792 6030 4809 6094
rect 4873 6030 4874 6094
rect 0 6008 4874 6030
rect 0 5944 105 6008
rect 169 5944 187 6008
rect 251 5944 269 6008
rect 333 5944 351 6008
rect 415 5944 433 6008
rect 497 5944 515 6008
rect 579 5944 597 6008
rect 661 5944 678 6008
rect 742 5944 759 6008
rect 823 5944 840 6008
rect 904 5944 921 6008
rect 985 5944 1002 6008
rect 1066 5944 1083 6008
rect 1147 5944 1164 6008
rect 1228 5944 1245 6008
rect 1309 5944 1326 6008
rect 1390 5944 1407 6008
rect 1471 5944 1488 6008
rect 1552 5944 1569 6008
rect 1633 5944 1650 6008
rect 1714 5944 1731 6008
rect 1795 5944 1812 6008
rect 1876 5944 1893 6008
rect 1957 5944 1974 6008
rect 2038 5944 2055 6008
rect 2119 5944 2136 6008
rect 2200 5944 2217 6008
rect 2281 5944 2298 6008
rect 2362 5944 2379 6008
rect 2443 5944 2460 6008
rect 2524 5944 2541 6008
rect 2605 5944 2622 6008
rect 2686 5944 2703 6008
rect 2767 5944 2784 6008
rect 2848 5944 2865 6008
rect 2929 5944 2946 6008
rect 3010 5944 3027 6008
rect 3091 5944 3108 6008
rect 3172 5944 3189 6008
rect 3253 5944 3270 6008
rect 3334 5944 3351 6008
rect 3415 5944 3432 6008
rect 3496 5944 3513 6008
rect 3577 5944 3594 6008
rect 3658 5944 3675 6008
rect 3739 5944 3756 6008
rect 3820 5944 3837 6008
rect 3901 5944 3918 6008
rect 3982 5944 3999 6008
rect 4063 5944 4080 6008
rect 4144 5944 4161 6008
rect 4225 5944 4242 6008
rect 4306 5944 4323 6008
rect 4387 5944 4404 6008
rect 4468 5944 4485 6008
rect 4549 5944 4566 6008
rect 4630 5944 4647 6008
rect 4711 5944 4728 6008
rect 4792 5944 4809 6008
rect 4873 5944 4874 6008
rect 0 5922 4874 5944
rect 0 5858 105 5922
rect 169 5858 187 5922
rect 251 5858 269 5922
rect 333 5858 351 5922
rect 415 5858 433 5922
rect 497 5858 515 5922
rect 579 5858 597 5922
rect 661 5858 678 5922
rect 742 5858 759 5922
rect 823 5858 840 5922
rect 904 5858 921 5922
rect 985 5858 1002 5922
rect 1066 5858 1083 5922
rect 1147 5858 1164 5922
rect 1228 5858 1245 5922
rect 1309 5858 1326 5922
rect 1390 5858 1407 5922
rect 1471 5858 1488 5922
rect 1552 5858 1569 5922
rect 1633 5858 1650 5922
rect 1714 5858 1731 5922
rect 1795 5858 1812 5922
rect 1876 5858 1893 5922
rect 1957 5858 1974 5922
rect 2038 5858 2055 5922
rect 2119 5858 2136 5922
rect 2200 5858 2217 5922
rect 2281 5858 2298 5922
rect 2362 5858 2379 5922
rect 2443 5858 2460 5922
rect 2524 5858 2541 5922
rect 2605 5858 2622 5922
rect 2686 5858 2703 5922
rect 2767 5858 2784 5922
rect 2848 5858 2865 5922
rect 2929 5858 2946 5922
rect 3010 5858 3027 5922
rect 3091 5858 3108 5922
rect 3172 5858 3189 5922
rect 3253 5858 3270 5922
rect 3334 5858 3351 5922
rect 3415 5858 3432 5922
rect 3496 5858 3513 5922
rect 3577 5858 3594 5922
rect 3658 5858 3675 5922
rect 3739 5858 3756 5922
rect 3820 5858 3837 5922
rect 3901 5858 3918 5922
rect 3982 5858 3999 5922
rect 4063 5858 4080 5922
rect 4144 5858 4161 5922
rect 4225 5858 4242 5922
rect 4306 5858 4323 5922
rect 4387 5858 4404 5922
rect 4468 5858 4485 5922
rect 4549 5858 4566 5922
rect 4630 5858 4647 5922
rect 4711 5858 4728 5922
rect 4792 5858 4809 5922
rect 4873 5858 4874 5922
rect 0 5836 4874 5858
rect 0 5772 105 5836
rect 169 5772 187 5836
rect 251 5772 269 5836
rect 333 5772 351 5836
rect 415 5772 433 5836
rect 497 5772 515 5836
rect 579 5772 597 5836
rect 661 5772 678 5836
rect 742 5772 759 5836
rect 823 5772 840 5836
rect 904 5772 921 5836
rect 985 5772 1002 5836
rect 1066 5772 1083 5836
rect 1147 5772 1164 5836
rect 1228 5772 1245 5836
rect 1309 5772 1326 5836
rect 1390 5772 1407 5836
rect 1471 5772 1488 5836
rect 1552 5772 1569 5836
rect 1633 5772 1650 5836
rect 1714 5772 1731 5836
rect 1795 5772 1812 5836
rect 1876 5772 1893 5836
rect 1957 5772 1974 5836
rect 2038 5772 2055 5836
rect 2119 5772 2136 5836
rect 2200 5772 2217 5836
rect 2281 5772 2298 5836
rect 2362 5772 2379 5836
rect 2443 5772 2460 5836
rect 2524 5772 2541 5836
rect 2605 5772 2622 5836
rect 2686 5772 2703 5836
rect 2767 5772 2784 5836
rect 2848 5772 2865 5836
rect 2929 5772 2946 5836
rect 3010 5772 3027 5836
rect 3091 5772 3108 5836
rect 3172 5772 3189 5836
rect 3253 5772 3270 5836
rect 3334 5772 3351 5836
rect 3415 5772 3432 5836
rect 3496 5772 3513 5836
rect 3577 5772 3594 5836
rect 3658 5772 3675 5836
rect 3739 5772 3756 5836
rect 3820 5772 3837 5836
rect 3901 5772 3918 5836
rect 3982 5772 3999 5836
rect 4063 5772 4080 5836
rect 4144 5772 4161 5836
rect 4225 5772 4242 5836
rect 4306 5772 4323 5836
rect 4387 5772 4404 5836
rect 4468 5772 4485 5836
rect 4549 5772 4566 5836
rect 4630 5772 4647 5836
rect 4711 5772 4728 5836
rect 4792 5772 4809 5836
rect 4873 5772 4874 5836
rect 0 5750 4874 5772
rect 0 5686 105 5750
rect 169 5686 187 5750
rect 251 5686 269 5750
rect 333 5686 351 5750
rect 415 5686 433 5750
rect 497 5686 515 5750
rect 579 5686 597 5750
rect 661 5686 678 5750
rect 742 5686 759 5750
rect 823 5686 840 5750
rect 904 5686 921 5750
rect 985 5686 1002 5750
rect 1066 5686 1083 5750
rect 1147 5686 1164 5750
rect 1228 5686 1245 5750
rect 1309 5686 1326 5750
rect 1390 5686 1407 5750
rect 1471 5686 1488 5750
rect 1552 5686 1569 5750
rect 1633 5686 1650 5750
rect 1714 5686 1731 5750
rect 1795 5686 1812 5750
rect 1876 5686 1893 5750
rect 1957 5686 1974 5750
rect 2038 5686 2055 5750
rect 2119 5686 2136 5750
rect 2200 5686 2217 5750
rect 2281 5686 2298 5750
rect 2362 5686 2379 5750
rect 2443 5686 2460 5750
rect 2524 5686 2541 5750
rect 2605 5686 2622 5750
rect 2686 5686 2703 5750
rect 2767 5686 2784 5750
rect 2848 5686 2865 5750
rect 2929 5686 2946 5750
rect 3010 5686 3027 5750
rect 3091 5686 3108 5750
rect 3172 5686 3189 5750
rect 3253 5686 3270 5750
rect 3334 5686 3351 5750
rect 3415 5686 3432 5750
rect 3496 5686 3513 5750
rect 3577 5686 3594 5750
rect 3658 5686 3675 5750
rect 3739 5686 3756 5750
rect 3820 5686 3837 5750
rect 3901 5686 3918 5750
rect 3982 5686 3999 5750
rect 4063 5686 4080 5750
rect 4144 5686 4161 5750
rect 4225 5686 4242 5750
rect 4306 5686 4323 5750
rect 4387 5686 4404 5750
rect 4468 5686 4485 5750
rect 4549 5686 4566 5750
rect 4630 5686 4647 5750
rect 4711 5686 4728 5750
rect 4792 5686 4809 5750
rect 4873 5686 4874 5750
rect 0 5664 4874 5686
rect 0 5600 105 5664
rect 169 5600 187 5664
rect 251 5600 269 5664
rect 333 5600 351 5664
rect 415 5600 433 5664
rect 497 5600 515 5664
rect 579 5600 597 5664
rect 661 5600 678 5664
rect 742 5600 759 5664
rect 823 5600 840 5664
rect 904 5600 921 5664
rect 985 5600 1002 5664
rect 1066 5600 1083 5664
rect 1147 5600 1164 5664
rect 1228 5600 1245 5664
rect 1309 5600 1326 5664
rect 1390 5600 1407 5664
rect 1471 5600 1488 5664
rect 1552 5600 1569 5664
rect 1633 5600 1650 5664
rect 1714 5600 1731 5664
rect 1795 5600 1812 5664
rect 1876 5600 1893 5664
rect 1957 5600 1974 5664
rect 2038 5600 2055 5664
rect 2119 5600 2136 5664
rect 2200 5600 2217 5664
rect 2281 5600 2298 5664
rect 2362 5600 2379 5664
rect 2443 5600 2460 5664
rect 2524 5600 2541 5664
rect 2605 5600 2622 5664
rect 2686 5600 2703 5664
rect 2767 5600 2784 5664
rect 2848 5600 2865 5664
rect 2929 5600 2946 5664
rect 3010 5600 3027 5664
rect 3091 5600 3108 5664
rect 3172 5600 3189 5664
rect 3253 5600 3270 5664
rect 3334 5600 3351 5664
rect 3415 5600 3432 5664
rect 3496 5600 3513 5664
rect 3577 5600 3594 5664
rect 3658 5600 3675 5664
rect 3739 5600 3756 5664
rect 3820 5600 3837 5664
rect 3901 5600 3918 5664
rect 3982 5600 3999 5664
rect 4063 5600 4080 5664
rect 4144 5600 4161 5664
rect 4225 5600 4242 5664
rect 4306 5600 4323 5664
rect 4387 5600 4404 5664
rect 4468 5600 4485 5664
rect 4549 5600 4566 5664
rect 4630 5600 4647 5664
rect 4711 5600 4728 5664
rect 4792 5600 4809 5664
rect 4873 5600 4874 5664
rect 0 5578 4874 5600
rect 0 5514 105 5578
rect 169 5514 187 5578
rect 251 5514 269 5578
rect 333 5514 351 5578
rect 415 5514 433 5578
rect 497 5514 515 5578
rect 579 5514 597 5578
rect 661 5514 678 5578
rect 742 5514 759 5578
rect 823 5514 840 5578
rect 904 5514 921 5578
rect 985 5514 1002 5578
rect 1066 5514 1083 5578
rect 1147 5514 1164 5578
rect 1228 5514 1245 5578
rect 1309 5514 1326 5578
rect 1390 5514 1407 5578
rect 1471 5514 1488 5578
rect 1552 5514 1569 5578
rect 1633 5514 1650 5578
rect 1714 5514 1731 5578
rect 1795 5514 1812 5578
rect 1876 5514 1893 5578
rect 1957 5514 1974 5578
rect 2038 5514 2055 5578
rect 2119 5514 2136 5578
rect 2200 5514 2217 5578
rect 2281 5514 2298 5578
rect 2362 5514 2379 5578
rect 2443 5514 2460 5578
rect 2524 5514 2541 5578
rect 2605 5514 2622 5578
rect 2686 5514 2703 5578
rect 2767 5514 2784 5578
rect 2848 5514 2865 5578
rect 2929 5514 2946 5578
rect 3010 5514 3027 5578
rect 3091 5514 3108 5578
rect 3172 5514 3189 5578
rect 3253 5514 3270 5578
rect 3334 5514 3351 5578
rect 3415 5514 3432 5578
rect 3496 5514 3513 5578
rect 3577 5514 3594 5578
rect 3658 5514 3675 5578
rect 3739 5514 3756 5578
rect 3820 5514 3837 5578
rect 3901 5514 3918 5578
rect 3982 5514 3999 5578
rect 4063 5514 4080 5578
rect 4144 5514 4161 5578
rect 4225 5514 4242 5578
rect 4306 5514 4323 5578
rect 4387 5514 4404 5578
rect 4468 5514 4485 5578
rect 4549 5514 4566 5578
rect 4630 5514 4647 5578
rect 4711 5514 4728 5578
rect 4792 5514 4809 5578
rect 4873 5514 4874 5578
rect 0 5492 4874 5514
rect 0 5428 105 5492
rect 169 5428 187 5492
rect 251 5428 269 5492
rect 333 5428 351 5492
rect 415 5428 433 5492
rect 497 5428 515 5492
rect 579 5428 597 5492
rect 661 5428 678 5492
rect 742 5428 759 5492
rect 823 5428 840 5492
rect 904 5428 921 5492
rect 985 5428 1002 5492
rect 1066 5428 1083 5492
rect 1147 5428 1164 5492
rect 1228 5428 1245 5492
rect 1309 5428 1326 5492
rect 1390 5428 1407 5492
rect 1471 5428 1488 5492
rect 1552 5428 1569 5492
rect 1633 5428 1650 5492
rect 1714 5428 1731 5492
rect 1795 5428 1812 5492
rect 1876 5428 1893 5492
rect 1957 5428 1974 5492
rect 2038 5428 2055 5492
rect 2119 5428 2136 5492
rect 2200 5428 2217 5492
rect 2281 5428 2298 5492
rect 2362 5428 2379 5492
rect 2443 5428 2460 5492
rect 2524 5428 2541 5492
rect 2605 5428 2622 5492
rect 2686 5428 2703 5492
rect 2767 5428 2784 5492
rect 2848 5428 2865 5492
rect 2929 5428 2946 5492
rect 3010 5428 3027 5492
rect 3091 5428 3108 5492
rect 3172 5428 3189 5492
rect 3253 5428 3270 5492
rect 3334 5428 3351 5492
rect 3415 5428 3432 5492
rect 3496 5428 3513 5492
rect 3577 5428 3594 5492
rect 3658 5428 3675 5492
rect 3739 5428 3756 5492
rect 3820 5428 3837 5492
rect 3901 5428 3918 5492
rect 3982 5428 3999 5492
rect 4063 5428 4080 5492
rect 4144 5428 4161 5492
rect 4225 5428 4242 5492
rect 4306 5428 4323 5492
rect 4387 5428 4404 5492
rect 4468 5428 4485 5492
rect 4549 5428 4566 5492
rect 4630 5428 4647 5492
rect 4711 5428 4728 5492
rect 4792 5428 4809 5492
rect 4873 5428 4874 5492
rect 0 5406 4874 5428
rect 0 5342 105 5406
rect 169 5342 187 5406
rect 251 5342 269 5406
rect 333 5342 351 5406
rect 415 5342 433 5406
rect 497 5342 515 5406
rect 579 5342 597 5406
rect 661 5342 678 5406
rect 742 5342 759 5406
rect 823 5342 840 5406
rect 904 5342 921 5406
rect 985 5342 1002 5406
rect 1066 5342 1083 5406
rect 1147 5342 1164 5406
rect 1228 5342 1245 5406
rect 1309 5342 1326 5406
rect 1390 5342 1407 5406
rect 1471 5342 1488 5406
rect 1552 5342 1569 5406
rect 1633 5342 1650 5406
rect 1714 5342 1731 5406
rect 1795 5342 1812 5406
rect 1876 5342 1893 5406
rect 1957 5342 1974 5406
rect 2038 5342 2055 5406
rect 2119 5342 2136 5406
rect 2200 5342 2217 5406
rect 2281 5342 2298 5406
rect 2362 5342 2379 5406
rect 2443 5342 2460 5406
rect 2524 5342 2541 5406
rect 2605 5342 2622 5406
rect 2686 5342 2703 5406
rect 2767 5342 2784 5406
rect 2848 5342 2865 5406
rect 2929 5342 2946 5406
rect 3010 5342 3027 5406
rect 3091 5342 3108 5406
rect 3172 5342 3189 5406
rect 3253 5342 3270 5406
rect 3334 5342 3351 5406
rect 3415 5342 3432 5406
rect 3496 5342 3513 5406
rect 3577 5342 3594 5406
rect 3658 5342 3675 5406
rect 3739 5342 3756 5406
rect 3820 5342 3837 5406
rect 3901 5342 3918 5406
rect 3982 5342 3999 5406
rect 4063 5342 4080 5406
rect 4144 5342 4161 5406
rect 4225 5342 4242 5406
rect 4306 5342 4323 5406
rect 4387 5342 4404 5406
rect 4468 5342 4485 5406
rect 4549 5342 4566 5406
rect 4630 5342 4647 5406
rect 4711 5342 4728 5406
rect 4792 5342 4809 5406
rect 4873 5342 4874 5406
rect 0 5320 4874 5342
rect 0 5256 105 5320
rect 169 5256 187 5320
rect 251 5256 269 5320
rect 333 5256 351 5320
rect 415 5256 433 5320
rect 497 5256 515 5320
rect 579 5256 597 5320
rect 661 5256 678 5320
rect 742 5256 759 5320
rect 823 5256 840 5320
rect 904 5256 921 5320
rect 985 5256 1002 5320
rect 1066 5256 1083 5320
rect 1147 5256 1164 5320
rect 1228 5256 1245 5320
rect 1309 5256 1326 5320
rect 1390 5256 1407 5320
rect 1471 5256 1488 5320
rect 1552 5256 1569 5320
rect 1633 5256 1650 5320
rect 1714 5256 1731 5320
rect 1795 5256 1812 5320
rect 1876 5256 1893 5320
rect 1957 5256 1974 5320
rect 2038 5256 2055 5320
rect 2119 5256 2136 5320
rect 2200 5256 2217 5320
rect 2281 5256 2298 5320
rect 2362 5256 2379 5320
rect 2443 5256 2460 5320
rect 2524 5256 2541 5320
rect 2605 5256 2622 5320
rect 2686 5256 2703 5320
rect 2767 5256 2784 5320
rect 2848 5256 2865 5320
rect 2929 5256 2946 5320
rect 3010 5256 3027 5320
rect 3091 5256 3108 5320
rect 3172 5256 3189 5320
rect 3253 5256 3270 5320
rect 3334 5256 3351 5320
rect 3415 5256 3432 5320
rect 3496 5256 3513 5320
rect 3577 5256 3594 5320
rect 3658 5256 3675 5320
rect 3739 5256 3756 5320
rect 3820 5256 3837 5320
rect 3901 5256 3918 5320
rect 3982 5256 3999 5320
rect 4063 5256 4080 5320
rect 4144 5256 4161 5320
rect 4225 5256 4242 5320
rect 4306 5256 4323 5320
rect 4387 5256 4404 5320
rect 4468 5256 4485 5320
rect 4549 5256 4566 5320
rect 4630 5256 4647 5320
rect 4711 5256 4728 5320
rect 4792 5256 4809 5320
rect 4873 5256 4874 5320
rect 0 5234 4874 5256
rect 0 5170 105 5234
rect 169 5170 187 5234
rect 251 5170 269 5234
rect 333 5170 351 5234
rect 415 5170 433 5234
rect 497 5170 515 5234
rect 579 5170 597 5234
rect 661 5170 678 5234
rect 742 5170 759 5234
rect 823 5170 840 5234
rect 904 5170 921 5234
rect 985 5170 1002 5234
rect 1066 5170 1083 5234
rect 1147 5170 1164 5234
rect 1228 5170 1245 5234
rect 1309 5170 1326 5234
rect 1390 5170 1407 5234
rect 1471 5170 1488 5234
rect 1552 5170 1569 5234
rect 1633 5170 1650 5234
rect 1714 5170 1731 5234
rect 1795 5170 1812 5234
rect 1876 5170 1893 5234
rect 1957 5170 1974 5234
rect 2038 5170 2055 5234
rect 2119 5170 2136 5234
rect 2200 5170 2217 5234
rect 2281 5170 2298 5234
rect 2362 5170 2379 5234
rect 2443 5170 2460 5234
rect 2524 5170 2541 5234
rect 2605 5170 2622 5234
rect 2686 5170 2703 5234
rect 2767 5170 2784 5234
rect 2848 5170 2865 5234
rect 2929 5170 2946 5234
rect 3010 5170 3027 5234
rect 3091 5170 3108 5234
rect 3172 5170 3189 5234
rect 3253 5170 3270 5234
rect 3334 5170 3351 5234
rect 3415 5170 3432 5234
rect 3496 5170 3513 5234
rect 3577 5170 3594 5234
rect 3658 5170 3675 5234
rect 3739 5170 3756 5234
rect 3820 5170 3837 5234
rect 3901 5170 3918 5234
rect 3982 5170 3999 5234
rect 4063 5170 4080 5234
rect 4144 5170 4161 5234
rect 4225 5170 4242 5234
rect 4306 5170 4323 5234
rect 4387 5170 4404 5234
rect 4468 5170 4485 5234
rect 4549 5170 4566 5234
rect 4630 5170 4647 5234
rect 4711 5170 4728 5234
rect 4792 5170 4809 5234
rect 4873 5170 4874 5234
rect 0 5167 4874 5170
rect 10083 6094 15000 6097
rect 10083 6030 10084 6094
rect 10148 6030 10166 6094
rect 10230 6030 10248 6094
rect 10312 6030 10330 6094
rect 10394 6030 10412 6094
rect 10476 6030 10494 6094
rect 10558 6030 10576 6094
rect 10640 6030 10657 6094
rect 10721 6030 10738 6094
rect 10802 6030 10819 6094
rect 10883 6030 10900 6094
rect 10964 6030 10981 6094
rect 11045 6030 11062 6094
rect 11126 6030 11143 6094
rect 11207 6030 11224 6094
rect 11288 6030 11305 6094
rect 11369 6030 11386 6094
rect 11450 6030 11467 6094
rect 11531 6030 11548 6094
rect 11612 6030 11629 6094
rect 11693 6030 11710 6094
rect 11774 6030 11791 6094
rect 11855 6030 11872 6094
rect 11936 6030 11953 6094
rect 12017 6030 12034 6094
rect 12098 6030 12115 6094
rect 12179 6030 12196 6094
rect 12260 6030 12277 6094
rect 12341 6030 12358 6094
rect 12422 6030 12439 6094
rect 12503 6030 12520 6094
rect 12584 6030 12601 6094
rect 12665 6030 12682 6094
rect 12746 6030 12763 6094
rect 12827 6030 12844 6094
rect 12908 6030 12925 6094
rect 12989 6030 13006 6094
rect 13070 6030 13087 6094
rect 13151 6030 13168 6094
rect 13232 6030 13249 6094
rect 13313 6030 13330 6094
rect 13394 6030 13411 6094
rect 13475 6030 13492 6094
rect 13556 6030 13573 6094
rect 13637 6030 13654 6094
rect 13718 6030 13735 6094
rect 13799 6030 13816 6094
rect 13880 6030 13897 6094
rect 13961 6030 13978 6094
rect 14042 6030 14059 6094
rect 14123 6030 14140 6094
rect 14204 6030 14221 6094
rect 14285 6030 14302 6094
rect 14366 6030 14383 6094
rect 14447 6030 14464 6094
rect 14528 6030 14545 6094
rect 14609 6030 14626 6094
rect 14690 6030 14707 6094
rect 14771 6030 14788 6094
rect 14852 6030 15000 6094
rect 10083 6008 15000 6030
rect 10083 5944 10084 6008
rect 10148 5944 10166 6008
rect 10230 5944 10248 6008
rect 10312 5944 10330 6008
rect 10394 5944 10412 6008
rect 10476 5944 10494 6008
rect 10558 5944 10576 6008
rect 10640 5944 10657 6008
rect 10721 5944 10738 6008
rect 10802 5944 10819 6008
rect 10883 5944 10900 6008
rect 10964 5944 10981 6008
rect 11045 5944 11062 6008
rect 11126 5944 11143 6008
rect 11207 5944 11224 6008
rect 11288 5944 11305 6008
rect 11369 5944 11386 6008
rect 11450 5944 11467 6008
rect 11531 5944 11548 6008
rect 11612 5944 11629 6008
rect 11693 5944 11710 6008
rect 11774 5944 11791 6008
rect 11855 5944 11872 6008
rect 11936 5944 11953 6008
rect 12017 5944 12034 6008
rect 12098 5944 12115 6008
rect 12179 5944 12196 6008
rect 12260 5944 12277 6008
rect 12341 5944 12358 6008
rect 12422 5944 12439 6008
rect 12503 5944 12520 6008
rect 12584 5944 12601 6008
rect 12665 5944 12682 6008
rect 12746 5944 12763 6008
rect 12827 5944 12844 6008
rect 12908 5944 12925 6008
rect 12989 5944 13006 6008
rect 13070 5944 13087 6008
rect 13151 5944 13168 6008
rect 13232 5944 13249 6008
rect 13313 5944 13330 6008
rect 13394 5944 13411 6008
rect 13475 5944 13492 6008
rect 13556 5944 13573 6008
rect 13637 5944 13654 6008
rect 13718 5944 13735 6008
rect 13799 5944 13816 6008
rect 13880 5944 13897 6008
rect 13961 5944 13978 6008
rect 14042 5944 14059 6008
rect 14123 5944 14140 6008
rect 14204 5944 14221 6008
rect 14285 5944 14302 6008
rect 14366 5944 14383 6008
rect 14447 5944 14464 6008
rect 14528 5944 14545 6008
rect 14609 5944 14626 6008
rect 14690 5944 14707 6008
rect 14771 5944 14788 6008
rect 14852 5944 15000 6008
rect 10083 5922 15000 5944
rect 10083 5858 10084 5922
rect 10148 5858 10166 5922
rect 10230 5858 10248 5922
rect 10312 5858 10330 5922
rect 10394 5858 10412 5922
rect 10476 5858 10494 5922
rect 10558 5858 10576 5922
rect 10640 5858 10657 5922
rect 10721 5858 10738 5922
rect 10802 5858 10819 5922
rect 10883 5858 10900 5922
rect 10964 5858 10981 5922
rect 11045 5858 11062 5922
rect 11126 5858 11143 5922
rect 11207 5858 11224 5922
rect 11288 5858 11305 5922
rect 11369 5858 11386 5922
rect 11450 5858 11467 5922
rect 11531 5858 11548 5922
rect 11612 5858 11629 5922
rect 11693 5858 11710 5922
rect 11774 5858 11791 5922
rect 11855 5858 11872 5922
rect 11936 5858 11953 5922
rect 12017 5858 12034 5922
rect 12098 5858 12115 5922
rect 12179 5858 12196 5922
rect 12260 5858 12277 5922
rect 12341 5858 12358 5922
rect 12422 5858 12439 5922
rect 12503 5858 12520 5922
rect 12584 5858 12601 5922
rect 12665 5858 12682 5922
rect 12746 5858 12763 5922
rect 12827 5858 12844 5922
rect 12908 5858 12925 5922
rect 12989 5858 13006 5922
rect 13070 5858 13087 5922
rect 13151 5858 13168 5922
rect 13232 5858 13249 5922
rect 13313 5858 13330 5922
rect 13394 5858 13411 5922
rect 13475 5858 13492 5922
rect 13556 5858 13573 5922
rect 13637 5858 13654 5922
rect 13718 5858 13735 5922
rect 13799 5858 13816 5922
rect 13880 5858 13897 5922
rect 13961 5858 13978 5922
rect 14042 5858 14059 5922
rect 14123 5858 14140 5922
rect 14204 5858 14221 5922
rect 14285 5858 14302 5922
rect 14366 5858 14383 5922
rect 14447 5858 14464 5922
rect 14528 5858 14545 5922
rect 14609 5858 14626 5922
rect 14690 5858 14707 5922
rect 14771 5858 14788 5922
rect 14852 5858 15000 5922
rect 10083 5836 15000 5858
rect 10083 5772 10084 5836
rect 10148 5772 10166 5836
rect 10230 5772 10248 5836
rect 10312 5772 10330 5836
rect 10394 5772 10412 5836
rect 10476 5772 10494 5836
rect 10558 5772 10576 5836
rect 10640 5772 10657 5836
rect 10721 5772 10738 5836
rect 10802 5772 10819 5836
rect 10883 5772 10900 5836
rect 10964 5772 10981 5836
rect 11045 5772 11062 5836
rect 11126 5772 11143 5836
rect 11207 5772 11224 5836
rect 11288 5772 11305 5836
rect 11369 5772 11386 5836
rect 11450 5772 11467 5836
rect 11531 5772 11548 5836
rect 11612 5772 11629 5836
rect 11693 5772 11710 5836
rect 11774 5772 11791 5836
rect 11855 5772 11872 5836
rect 11936 5772 11953 5836
rect 12017 5772 12034 5836
rect 12098 5772 12115 5836
rect 12179 5772 12196 5836
rect 12260 5772 12277 5836
rect 12341 5772 12358 5836
rect 12422 5772 12439 5836
rect 12503 5772 12520 5836
rect 12584 5772 12601 5836
rect 12665 5772 12682 5836
rect 12746 5772 12763 5836
rect 12827 5772 12844 5836
rect 12908 5772 12925 5836
rect 12989 5772 13006 5836
rect 13070 5772 13087 5836
rect 13151 5772 13168 5836
rect 13232 5772 13249 5836
rect 13313 5772 13330 5836
rect 13394 5772 13411 5836
rect 13475 5772 13492 5836
rect 13556 5772 13573 5836
rect 13637 5772 13654 5836
rect 13718 5772 13735 5836
rect 13799 5772 13816 5836
rect 13880 5772 13897 5836
rect 13961 5772 13978 5836
rect 14042 5772 14059 5836
rect 14123 5772 14140 5836
rect 14204 5772 14221 5836
rect 14285 5772 14302 5836
rect 14366 5772 14383 5836
rect 14447 5772 14464 5836
rect 14528 5772 14545 5836
rect 14609 5772 14626 5836
rect 14690 5772 14707 5836
rect 14771 5772 14788 5836
rect 14852 5772 15000 5836
rect 10083 5750 15000 5772
rect 10083 5686 10084 5750
rect 10148 5686 10166 5750
rect 10230 5686 10248 5750
rect 10312 5686 10330 5750
rect 10394 5686 10412 5750
rect 10476 5686 10494 5750
rect 10558 5686 10576 5750
rect 10640 5686 10657 5750
rect 10721 5686 10738 5750
rect 10802 5686 10819 5750
rect 10883 5686 10900 5750
rect 10964 5686 10981 5750
rect 11045 5686 11062 5750
rect 11126 5686 11143 5750
rect 11207 5686 11224 5750
rect 11288 5686 11305 5750
rect 11369 5686 11386 5750
rect 11450 5686 11467 5750
rect 11531 5686 11548 5750
rect 11612 5686 11629 5750
rect 11693 5686 11710 5750
rect 11774 5686 11791 5750
rect 11855 5686 11872 5750
rect 11936 5686 11953 5750
rect 12017 5686 12034 5750
rect 12098 5686 12115 5750
rect 12179 5686 12196 5750
rect 12260 5686 12277 5750
rect 12341 5686 12358 5750
rect 12422 5686 12439 5750
rect 12503 5686 12520 5750
rect 12584 5686 12601 5750
rect 12665 5686 12682 5750
rect 12746 5686 12763 5750
rect 12827 5686 12844 5750
rect 12908 5686 12925 5750
rect 12989 5686 13006 5750
rect 13070 5686 13087 5750
rect 13151 5686 13168 5750
rect 13232 5686 13249 5750
rect 13313 5686 13330 5750
rect 13394 5686 13411 5750
rect 13475 5686 13492 5750
rect 13556 5686 13573 5750
rect 13637 5686 13654 5750
rect 13718 5686 13735 5750
rect 13799 5686 13816 5750
rect 13880 5686 13897 5750
rect 13961 5686 13978 5750
rect 14042 5686 14059 5750
rect 14123 5686 14140 5750
rect 14204 5686 14221 5750
rect 14285 5686 14302 5750
rect 14366 5686 14383 5750
rect 14447 5686 14464 5750
rect 14528 5686 14545 5750
rect 14609 5686 14626 5750
rect 14690 5686 14707 5750
rect 14771 5686 14788 5750
rect 14852 5686 15000 5750
rect 10083 5664 15000 5686
rect 10083 5600 10084 5664
rect 10148 5600 10166 5664
rect 10230 5600 10248 5664
rect 10312 5600 10330 5664
rect 10394 5600 10412 5664
rect 10476 5600 10494 5664
rect 10558 5600 10576 5664
rect 10640 5600 10657 5664
rect 10721 5600 10738 5664
rect 10802 5600 10819 5664
rect 10883 5600 10900 5664
rect 10964 5600 10981 5664
rect 11045 5600 11062 5664
rect 11126 5600 11143 5664
rect 11207 5600 11224 5664
rect 11288 5600 11305 5664
rect 11369 5600 11386 5664
rect 11450 5600 11467 5664
rect 11531 5600 11548 5664
rect 11612 5600 11629 5664
rect 11693 5600 11710 5664
rect 11774 5600 11791 5664
rect 11855 5600 11872 5664
rect 11936 5600 11953 5664
rect 12017 5600 12034 5664
rect 12098 5600 12115 5664
rect 12179 5600 12196 5664
rect 12260 5600 12277 5664
rect 12341 5600 12358 5664
rect 12422 5600 12439 5664
rect 12503 5600 12520 5664
rect 12584 5600 12601 5664
rect 12665 5600 12682 5664
rect 12746 5600 12763 5664
rect 12827 5600 12844 5664
rect 12908 5600 12925 5664
rect 12989 5600 13006 5664
rect 13070 5600 13087 5664
rect 13151 5600 13168 5664
rect 13232 5600 13249 5664
rect 13313 5600 13330 5664
rect 13394 5600 13411 5664
rect 13475 5600 13492 5664
rect 13556 5600 13573 5664
rect 13637 5600 13654 5664
rect 13718 5600 13735 5664
rect 13799 5600 13816 5664
rect 13880 5600 13897 5664
rect 13961 5600 13978 5664
rect 14042 5600 14059 5664
rect 14123 5600 14140 5664
rect 14204 5600 14221 5664
rect 14285 5600 14302 5664
rect 14366 5600 14383 5664
rect 14447 5600 14464 5664
rect 14528 5600 14545 5664
rect 14609 5600 14626 5664
rect 14690 5600 14707 5664
rect 14771 5600 14788 5664
rect 14852 5600 15000 5664
rect 10083 5578 15000 5600
rect 10083 5514 10084 5578
rect 10148 5514 10166 5578
rect 10230 5514 10248 5578
rect 10312 5514 10330 5578
rect 10394 5514 10412 5578
rect 10476 5514 10494 5578
rect 10558 5514 10576 5578
rect 10640 5514 10657 5578
rect 10721 5514 10738 5578
rect 10802 5514 10819 5578
rect 10883 5514 10900 5578
rect 10964 5514 10981 5578
rect 11045 5514 11062 5578
rect 11126 5514 11143 5578
rect 11207 5514 11224 5578
rect 11288 5514 11305 5578
rect 11369 5514 11386 5578
rect 11450 5514 11467 5578
rect 11531 5514 11548 5578
rect 11612 5514 11629 5578
rect 11693 5514 11710 5578
rect 11774 5514 11791 5578
rect 11855 5514 11872 5578
rect 11936 5514 11953 5578
rect 12017 5514 12034 5578
rect 12098 5514 12115 5578
rect 12179 5514 12196 5578
rect 12260 5514 12277 5578
rect 12341 5514 12358 5578
rect 12422 5514 12439 5578
rect 12503 5514 12520 5578
rect 12584 5514 12601 5578
rect 12665 5514 12682 5578
rect 12746 5514 12763 5578
rect 12827 5514 12844 5578
rect 12908 5514 12925 5578
rect 12989 5514 13006 5578
rect 13070 5514 13087 5578
rect 13151 5514 13168 5578
rect 13232 5514 13249 5578
rect 13313 5514 13330 5578
rect 13394 5514 13411 5578
rect 13475 5514 13492 5578
rect 13556 5514 13573 5578
rect 13637 5514 13654 5578
rect 13718 5514 13735 5578
rect 13799 5514 13816 5578
rect 13880 5514 13897 5578
rect 13961 5514 13978 5578
rect 14042 5514 14059 5578
rect 14123 5514 14140 5578
rect 14204 5514 14221 5578
rect 14285 5514 14302 5578
rect 14366 5514 14383 5578
rect 14447 5514 14464 5578
rect 14528 5514 14545 5578
rect 14609 5514 14626 5578
rect 14690 5514 14707 5578
rect 14771 5514 14788 5578
rect 14852 5514 15000 5578
rect 10083 5492 15000 5514
rect 10083 5428 10084 5492
rect 10148 5428 10166 5492
rect 10230 5428 10248 5492
rect 10312 5428 10330 5492
rect 10394 5428 10412 5492
rect 10476 5428 10494 5492
rect 10558 5428 10576 5492
rect 10640 5428 10657 5492
rect 10721 5428 10738 5492
rect 10802 5428 10819 5492
rect 10883 5428 10900 5492
rect 10964 5428 10981 5492
rect 11045 5428 11062 5492
rect 11126 5428 11143 5492
rect 11207 5428 11224 5492
rect 11288 5428 11305 5492
rect 11369 5428 11386 5492
rect 11450 5428 11467 5492
rect 11531 5428 11548 5492
rect 11612 5428 11629 5492
rect 11693 5428 11710 5492
rect 11774 5428 11791 5492
rect 11855 5428 11872 5492
rect 11936 5428 11953 5492
rect 12017 5428 12034 5492
rect 12098 5428 12115 5492
rect 12179 5428 12196 5492
rect 12260 5428 12277 5492
rect 12341 5428 12358 5492
rect 12422 5428 12439 5492
rect 12503 5428 12520 5492
rect 12584 5428 12601 5492
rect 12665 5428 12682 5492
rect 12746 5428 12763 5492
rect 12827 5428 12844 5492
rect 12908 5428 12925 5492
rect 12989 5428 13006 5492
rect 13070 5428 13087 5492
rect 13151 5428 13168 5492
rect 13232 5428 13249 5492
rect 13313 5428 13330 5492
rect 13394 5428 13411 5492
rect 13475 5428 13492 5492
rect 13556 5428 13573 5492
rect 13637 5428 13654 5492
rect 13718 5428 13735 5492
rect 13799 5428 13816 5492
rect 13880 5428 13897 5492
rect 13961 5428 13978 5492
rect 14042 5428 14059 5492
rect 14123 5428 14140 5492
rect 14204 5428 14221 5492
rect 14285 5428 14302 5492
rect 14366 5428 14383 5492
rect 14447 5428 14464 5492
rect 14528 5428 14545 5492
rect 14609 5428 14626 5492
rect 14690 5428 14707 5492
rect 14771 5428 14788 5492
rect 14852 5428 15000 5492
rect 10083 5406 15000 5428
rect 10083 5342 10084 5406
rect 10148 5342 10166 5406
rect 10230 5342 10248 5406
rect 10312 5342 10330 5406
rect 10394 5342 10412 5406
rect 10476 5342 10494 5406
rect 10558 5342 10576 5406
rect 10640 5342 10657 5406
rect 10721 5342 10738 5406
rect 10802 5342 10819 5406
rect 10883 5342 10900 5406
rect 10964 5342 10981 5406
rect 11045 5342 11062 5406
rect 11126 5342 11143 5406
rect 11207 5342 11224 5406
rect 11288 5342 11305 5406
rect 11369 5342 11386 5406
rect 11450 5342 11467 5406
rect 11531 5342 11548 5406
rect 11612 5342 11629 5406
rect 11693 5342 11710 5406
rect 11774 5342 11791 5406
rect 11855 5342 11872 5406
rect 11936 5342 11953 5406
rect 12017 5342 12034 5406
rect 12098 5342 12115 5406
rect 12179 5342 12196 5406
rect 12260 5342 12277 5406
rect 12341 5342 12358 5406
rect 12422 5342 12439 5406
rect 12503 5342 12520 5406
rect 12584 5342 12601 5406
rect 12665 5342 12682 5406
rect 12746 5342 12763 5406
rect 12827 5342 12844 5406
rect 12908 5342 12925 5406
rect 12989 5342 13006 5406
rect 13070 5342 13087 5406
rect 13151 5342 13168 5406
rect 13232 5342 13249 5406
rect 13313 5342 13330 5406
rect 13394 5342 13411 5406
rect 13475 5342 13492 5406
rect 13556 5342 13573 5406
rect 13637 5342 13654 5406
rect 13718 5342 13735 5406
rect 13799 5342 13816 5406
rect 13880 5342 13897 5406
rect 13961 5342 13978 5406
rect 14042 5342 14059 5406
rect 14123 5342 14140 5406
rect 14204 5342 14221 5406
rect 14285 5342 14302 5406
rect 14366 5342 14383 5406
rect 14447 5342 14464 5406
rect 14528 5342 14545 5406
rect 14609 5342 14626 5406
rect 14690 5342 14707 5406
rect 14771 5342 14788 5406
rect 14852 5342 15000 5406
rect 10083 5320 15000 5342
rect 10083 5256 10084 5320
rect 10148 5256 10166 5320
rect 10230 5256 10248 5320
rect 10312 5256 10330 5320
rect 10394 5256 10412 5320
rect 10476 5256 10494 5320
rect 10558 5256 10576 5320
rect 10640 5256 10657 5320
rect 10721 5256 10738 5320
rect 10802 5256 10819 5320
rect 10883 5256 10900 5320
rect 10964 5256 10981 5320
rect 11045 5256 11062 5320
rect 11126 5256 11143 5320
rect 11207 5256 11224 5320
rect 11288 5256 11305 5320
rect 11369 5256 11386 5320
rect 11450 5256 11467 5320
rect 11531 5256 11548 5320
rect 11612 5256 11629 5320
rect 11693 5256 11710 5320
rect 11774 5256 11791 5320
rect 11855 5256 11872 5320
rect 11936 5256 11953 5320
rect 12017 5256 12034 5320
rect 12098 5256 12115 5320
rect 12179 5256 12196 5320
rect 12260 5256 12277 5320
rect 12341 5256 12358 5320
rect 12422 5256 12439 5320
rect 12503 5256 12520 5320
rect 12584 5256 12601 5320
rect 12665 5256 12682 5320
rect 12746 5256 12763 5320
rect 12827 5256 12844 5320
rect 12908 5256 12925 5320
rect 12989 5256 13006 5320
rect 13070 5256 13087 5320
rect 13151 5256 13168 5320
rect 13232 5256 13249 5320
rect 13313 5256 13330 5320
rect 13394 5256 13411 5320
rect 13475 5256 13492 5320
rect 13556 5256 13573 5320
rect 13637 5256 13654 5320
rect 13718 5256 13735 5320
rect 13799 5256 13816 5320
rect 13880 5256 13897 5320
rect 13961 5256 13978 5320
rect 14042 5256 14059 5320
rect 14123 5256 14140 5320
rect 14204 5256 14221 5320
rect 14285 5256 14302 5320
rect 14366 5256 14383 5320
rect 14447 5256 14464 5320
rect 14528 5256 14545 5320
rect 14609 5256 14626 5320
rect 14690 5256 14707 5320
rect 14771 5256 14788 5320
rect 14852 5256 15000 5320
rect 10083 5234 15000 5256
rect 10083 5170 10084 5234
rect 10148 5170 10166 5234
rect 10230 5170 10248 5234
rect 10312 5170 10330 5234
rect 10394 5170 10412 5234
rect 10476 5170 10494 5234
rect 10558 5170 10576 5234
rect 10640 5170 10657 5234
rect 10721 5170 10738 5234
rect 10802 5170 10819 5234
rect 10883 5170 10900 5234
rect 10964 5170 10981 5234
rect 11045 5170 11062 5234
rect 11126 5170 11143 5234
rect 11207 5170 11224 5234
rect 11288 5170 11305 5234
rect 11369 5170 11386 5234
rect 11450 5170 11467 5234
rect 11531 5170 11548 5234
rect 11612 5170 11629 5234
rect 11693 5170 11710 5234
rect 11774 5170 11791 5234
rect 11855 5170 11872 5234
rect 11936 5170 11953 5234
rect 12017 5170 12034 5234
rect 12098 5170 12115 5234
rect 12179 5170 12196 5234
rect 12260 5170 12277 5234
rect 12341 5170 12358 5234
rect 12422 5170 12439 5234
rect 12503 5170 12520 5234
rect 12584 5170 12601 5234
rect 12665 5170 12682 5234
rect 12746 5170 12763 5234
rect 12827 5170 12844 5234
rect 12908 5170 12925 5234
rect 12989 5170 13006 5234
rect 13070 5170 13087 5234
rect 13151 5170 13168 5234
rect 13232 5170 13249 5234
rect 13313 5170 13330 5234
rect 13394 5170 13411 5234
rect 13475 5170 13492 5234
rect 13556 5170 13573 5234
rect 13637 5170 13654 5234
rect 13718 5170 13735 5234
rect 13799 5170 13816 5234
rect 13880 5170 13897 5234
rect 13961 5170 13978 5234
rect 14042 5170 14059 5234
rect 14123 5170 14140 5234
rect 14204 5170 14221 5234
rect 14285 5170 14302 5234
rect 14366 5170 14383 5234
rect 14447 5170 14464 5234
rect 14528 5170 14545 5234
rect 14609 5170 14626 5234
rect 14690 5170 14707 5234
rect 14771 5170 14788 5234
rect 14852 5170 15000 5234
rect 10083 5167 15000 5170
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 14746 14007 15000 18997
rect 0 12837 254 13687
rect 14746 12837 15000 13687
rect 0 11667 254 12517
rect 14746 11667 15000 12517
rect 0 9547 254 11347
rect 14746 9547 15000 11347
rect 0 8337 254 9227
rect 14746 8337 15000 9227
rect 0 7368 254 8017
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 14746 6397 15000 7047
rect 0 5187 254 6077
rect 14746 5187 15000 6077
rect 0 3977 254 4867
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 14746 1797 15000 2687
rect 0 427 254 1477
rect 14746 427 15000 1477
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1676037725
transform 1 0 0 0 1 549
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 28 nsew ground bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 16 nsew power bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 24 nsew power bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 29 nsew ground bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 40 nsew ground bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 44 nsew ground bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 56 nsew power bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 52 nsew ground bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 17 nsew power bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 12 nsew power bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 4 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 8 nsew power bidirectional
flabel metal5 s 14746 9547 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 30 nsew ground bidirectional
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 520 180 0 0 VDDIO
port 18 nsew power bidirectional
flabel metal5 s 14746 12837 15000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 25 nsew power bidirectional
flabel metal5 s 14746 7368 15000 8017 3 FreeSans 520 180 0 0 VSSA
port 31 nsew ground bidirectional
flabel metal5 s 14746 8337 15000 9227 3 FreeSans 520 180 0 0 VSSD
port 41 nsew ground bidirectional
flabel metal5 s 14746 5187 15000 6077 3 FreeSans 520 180 0 0 VSSIO
port 45 nsew ground bidirectional
flabel metal5 s 14746 6397 15000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 57 nsew power bidirectional
flabel metal5 s 14746 11667 15000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 53 nsew ground bidirectional
flabel metal5 s 14746 3977 15000 4867 3 FreeSans 520 180 0 0 VDDIO
port 19 nsew power bidirectional
flabel metal5 s 14807 3007 15000 3657 3 FreeSans 520 180 0 0 VDDA
port 13 nsew power bidirectional
flabel metal5 s 14746 1797 15000 2687 3 FreeSans 520 180 0 0 VCCD
port 5 nsew power bidirectional
flabel metal5 s 14746 427 15000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 46 nsew ground bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 47 nsew ground bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 20 nsew power bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 32 nsew ground bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 58 nsew power bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 48 nsew ground bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 54 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 34 nsew ground bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 14 nsew power bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 6 nsew power bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 10 nsew power bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 2 nsew signal bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 26 nsew power bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 42 nsew ground bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 35 nsew ground bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 0 nsew signal bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 21 nsew power bidirectional
flabel metal4 s 14746 3957 15000 4887 3 FreeSans 520 180 0 0 VDDIO
port 22 nsew power bidirectional
flabel metal4 s 14746 11281 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 36 nsew ground bidirectional
flabel metal4 s 14746 6377 15000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 59 nsew power bidirectional
flabel metal4 s 14746 5167 15000 6097 3 FreeSans 520 180 0 0 VSSIO
port 49 nsew ground bidirectional
flabel metal4 s 14746 11647 15000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 55 nsew ground bidirectional
flabel metal4 s 14746 9547 15000 9613 3 FreeSans 520 180 0 0 VSSA
port 37 nsew ground bidirectional
flabel metal4 s 14746 10329 15000 10565 3 FreeSans 520 180 0 0 VSSA
port 38 nsew ground bidirectional
flabel metal4 s 14807 2987 15000 3677 3 FreeSans 520 180 0 0 VDDA
port 15 nsew power bidirectional
flabel metal4 s 14746 1777 15000 2707 3 FreeSans 520 180 0 0 VCCD
port 7 nsew power bidirectional
flabel metal4 s 14746 407 15000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 11 nsew power bidirectional
flabel metal4 s 14746 9673 15000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 3 nsew signal bidirectional
flabel metal4 s 14746 12817 15000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 27 nsew power bidirectional
flabel metal4 s 14746 8317 15000 9247 3 FreeSans 520 180 0 0 VSSD
port 43 nsew ground bidirectional
flabel metal4 s 14746 7347 15000 8037 3 FreeSans 520 180 0 0 VSSA
port 39 nsew ground bidirectional
flabel metal4 s 14746 10625 15000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 1 nsew signal bidirectional
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 520 180 0 0 VDDIO
port 23 nsew power bidirectional
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 50 nsew ground bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 51 nsew ground bidirectional
flabel metal4 s 127 38321 127 38321 3 FreeSans 520 0 0 0 VSSIO
rlabel metal4 s 14746 10625 15000 11221 1 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 1 AMUXBUS_B
port 3 nsew signal bidirectional
rlabel metal4 s 14746 1777 15000 2707 1 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 1 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 1 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 1 VCCHIB
port 11 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 1 VCCHIB
port 11 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 1 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 1 VDDA
port 15 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 1 VDDA
port 15 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 1 VDDA
port 15 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 1 VDDIO
port 23 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 1 VDDIO
port 23 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 1 VDDIO
port 23 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 1 VDDIO
port 23 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 1 VDDIO
port 23 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 1 VDDIO
port 23 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 1 VDDIO
port 23 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 1 VDDIO_Q
port 27 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 1 VDDIO_Q
port 27 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 1 VDDIO_Q
port 27 nsew power bidirectional
rlabel metal4 s 0 9547 254 9613 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 1 VSSA
port 39 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 1 VSSA
port 39 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 1 VSSA
port 39 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 1 VSSA
port 39 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 1 VSSD
port 43 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 1 VSSD
port 43 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 1 VSSD
port 43 nsew ground bidirectional
rlabel metal3 s 99 5168 4879 6096 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal3 s 10078 5168 14858 6096 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 0 39984 254 40000 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 0 35186 2695 39984 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 0 35157 254 35186 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 0 5167 4874 6097 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 2719 39246 2851 39394 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 2726 39434 12265 39986 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 10083 5167 15000 6097 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 12136 39246 12268 39394 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 14746 39984 15000 40000 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 35186 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal4 s 12301 35186 15000 39984 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 6042 14840 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5956 14840 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5870 14840 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5784 14840 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5698 14840 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5612 14840 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5526 14840 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5440 14840 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5354 14840 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5268 14840 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14800 5182 14840 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39931 14838 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39850 14838 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39769 14838 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39688 14838 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39607 14838 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39526 14838 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39445 14838 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39364 14838 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39283 14838 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39202 14838 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39121 14838 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 39040 14838 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38959 14838 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38879 14838 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38799 14838 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38719 14838 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38639 14838 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38559 14838 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38479 14838 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38399 14838 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38319 14838 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38239 14838 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38159 14838 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 38079 14838 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37999 14838 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37919 14838 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37839 14838 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37759 14838 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37679 14838 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37599 14838 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37519 14838 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37439 14838 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37359 14838 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37279 14838 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37199 14838 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37119 14838 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 37039 14838 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36959 14838 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36879 14838 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36799 14838 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36719 14838 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36639 14838 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36559 14838 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36479 14838 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36399 14838 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36319 14838 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36239 14838 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36159 14838 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 36079 14838 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35999 14838 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35919 14838 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35839 14838 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35759 14838 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35679 14838 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35599 14838 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35519 14838 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35439 14838 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35359 14838 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35279 14838 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14798 35199 14838 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 6042 14759 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5956 14759 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5870 14759 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5784 14759 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5698 14759 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5612 14759 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5526 14759 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5440 14759 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5354 14759 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5268 14759 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14719 5182 14759 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39931 14758 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39850 14758 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39769 14758 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39688 14758 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39607 14758 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39526 14758 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39445 14758 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39364 14758 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39283 14758 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39202 14758 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39121 14758 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 39040 14758 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38959 14758 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38879 14758 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38799 14758 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38719 14758 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38639 14758 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38559 14758 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38479 14758 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38399 14758 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38319 14758 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38239 14758 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38159 14758 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 38079 14758 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37999 14758 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37919 14758 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37839 14758 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37759 14758 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37679 14758 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37599 14758 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37519 14758 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37439 14758 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37359 14758 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37279 14758 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37199 14758 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37119 14758 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 37039 14758 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36959 14758 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36879 14758 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36799 14758 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36719 14758 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36639 14758 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36559 14758 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36479 14758 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36399 14758 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36319 14758 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36239 14758 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36159 14758 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 36079 14758 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35999 14758 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35919 14758 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35839 14758 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35759 14758 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35679 14758 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35599 14758 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35519 14758 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35439 14758 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35359 14758 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35279 14758 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14718 35199 14758 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39931 14678 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39850 14678 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39769 14678 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39688 14678 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39607 14678 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39526 14678 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39445 14678 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39364 14678 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39283 14678 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39202 14678 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39121 14678 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 39040 14678 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38959 14678 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38879 14678 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38799 14678 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38719 14678 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38639 14678 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38559 14678 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38479 14678 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38399 14678 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38319 14678 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38239 14678 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38159 14678 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 38079 14678 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37999 14678 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37919 14678 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37839 14678 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37759 14678 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37679 14678 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37599 14678 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37519 14678 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37439 14678 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37359 14678 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37279 14678 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37199 14678 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37119 14678 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 37039 14678 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36959 14678 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36879 14678 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36799 14678 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36719 14678 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36639 14678 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36559 14678 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36479 14678 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36399 14678 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36319 14678 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36239 14678 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36159 14678 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 36079 14678 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35999 14678 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35919 14678 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35839 14678 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35759 14678 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35679 14678 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35599 14678 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35519 14678 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35439 14678 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35359 14678 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35279 14678 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 35199 14678 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 6042 14678 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5956 14678 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5870 14678 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5784 14678 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5698 14678 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5612 14678 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5526 14678 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5440 14678 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5354 14678 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5268 14678 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14638 5182 14678 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39931 14598 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39850 14598 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39769 14598 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39688 14598 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39607 14598 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39526 14598 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39445 14598 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39364 14598 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39283 14598 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39202 14598 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39121 14598 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 39040 14598 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38959 14598 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38879 14598 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38799 14598 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38719 14598 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38639 14598 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38559 14598 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38479 14598 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38399 14598 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38319 14598 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38239 14598 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38159 14598 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 38079 14598 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37999 14598 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37919 14598 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37839 14598 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37759 14598 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37679 14598 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37599 14598 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37519 14598 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37439 14598 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37359 14598 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37279 14598 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37199 14598 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37119 14598 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 37039 14598 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36959 14598 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36879 14598 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36799 14598 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36719 14598 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36639 14598 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36559 14598 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36479 14598 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36399 14598 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36319 14598 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36239 14598 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36159 14598 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 36079 14598 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35999 14598 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35919 14598 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35839 14598 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35759 14598 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35679 14598 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35599 14598 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35519 14598 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35439 14598 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35359 14598 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35279 14598 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14558 35199 14598 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 6042 14597 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5956 14597 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5870 14597 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5784 14597 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5698 14597 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5612 14597 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5526 14597 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5440 14597 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5354 14597 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5268 14597 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14557 5182 14597 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39931 14518 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39850 14518 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39769 14518 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39688 14518 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39607 14518 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39526 14518 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39445 14518 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39364 14518 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39283 14518 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39202 14518 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39121 14518 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 39040 14518 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38959 14518 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38879 14518 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38799 14518 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38719 14518 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38639 14518 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38559 14518 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38479 14518 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38399 14518 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38319 14518 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38239 14518 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38159 14518 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 38079 14518 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37999 14518 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37919 14518 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37839 14518 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37759 14518 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37679 14518 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37599 14518 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37519 14518 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37439 14518 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37359 14518 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37279 14518 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37199 14518 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37119 14518 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 37039 14518 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36959 14518 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36879 14518 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36799 14518 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36719 14518 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36639 14518 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36559 14518 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36479 14518 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36399 14518 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36319 14518 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36239 14518 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36159 14518 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 36079 14518 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35999 14518 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35919 14518 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35839 14518 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35759 14518 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35679 14518 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35599 14518 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35519 14518 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35439 14518 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35359 14518 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35279 14518 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14478 35199 14518 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 6042 14516 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5956 14516 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5870 14516 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5784 14516 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5698 14516 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5612 14516 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5526 14516 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5440 14516 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5354 14516 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5268 14516 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14476 5182 14516 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39931 14438 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39850 14438 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39769 14438 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39688 14438 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39607 14438 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39526 14438 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39445 14438 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39364 14438 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39283 14438 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39202 14438 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39121 14438 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 39040 14438 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38959 14438 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38879 14438 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38799 14438 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38719 14438 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38639 14438 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38559 14438 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38479 14438 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38399 14438 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38319 14438 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38239 14438 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38159 14438 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 38079 14438 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37999 14438 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37919 14438 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37839 14438 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37759 14438 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37679 14438 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37599 14438 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37519 14438 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37439 14438 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37359 14438 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37279 14438 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37199 14438 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37119 14438 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 37039 14438 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36959 14438 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36879 14438 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36799 14438 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36719 14438 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36639 14438 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36559 14438 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36479 14438 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36399 14438 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36319 14438 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36239 14438 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36159 14438 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 36079 14438 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35999 14438 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35919 14438 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35839 14438 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35759 14438 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35679 14438 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35599 14438 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35519 14438 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35439 14438 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35359 14438 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35279 14438 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14398 35199 14438 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 6042 14435 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5956 14435 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5870 14435 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5784 14435 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5698 14435 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5612 14435 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5526 14435 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5440 14435 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5354 14435 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5268 14435 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14395 5182 14435 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39931 14358 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39850 14358 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39769 14358 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39688 14358 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39607 14358 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39526 14358 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39445 14358 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39364 14358 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39283 14358 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39202 14358 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39121 14358 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 39040 14358 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38959 14358 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38879 14358 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38799 14358 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38719 14358 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38639 14358 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38559 14358 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38479 14358 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38399 14358 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38319 14358 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38239 14358 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38159 14358 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 38079 14358 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37999 14358 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37919 14358 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37839 14358 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37759 14358 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37679 14358 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37599 14358 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37519 14358 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37439 14358 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37359 14358 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37279 14358 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37199 14358 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37119 14358 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 37039 14358 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36959 14358 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36879 14358 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36799 14358 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36719 14358 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36639 14358 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36559 14358 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36479 14358 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36399 14358 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36319 14358 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36239 14358 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36159 14358 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 36079 14358 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35999 14358 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35919 14358 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35839 14358 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35759 14358 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35679 14358 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35599 14358 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35519 14358 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35439 14358 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35359 14358 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35279 14358 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14318 35199 14358 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 6042 14354 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5956 14354 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5870 14354 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5784 14354 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5698 14354 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5612 14354 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5526 14354 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5440 14354 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5354 14354 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5268 14354 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14314 5182 14354 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39931 14278 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39850 14278 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39769 14278 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39688 14278 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39607 14278 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39526 14278 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39445 14278 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39364 14278 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39283 14278 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39202 14278 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39121 14278 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 39040 14278 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38959 14278 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38879 14278 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38799 14278 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38719 14278 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38639 14278 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38559 14278 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38479 14278 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38399 14278 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38319 14278 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38239 14278 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38159 14278 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 38079 14278 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37999 14278 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37919 14278 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37839 14278 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37759 14278 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37679 14278 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37599 14278 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37519 14278 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37439 14278 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37359 14278 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37279 14278 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37199 14278 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37119 14278 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 37039 14278 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36959 14278 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36879 14278 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36799 14278 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36719 14278 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36639 14278 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36559 14278 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36479 14278 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36399 14278 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36319 14278 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36239 14278 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36159 14278 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 36079 14278 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35999 14278 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35919 14278 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35839 14278 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35759 14278 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35679 14278 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35599 14278 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35519 14278 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35439 14278 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35359 14278 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35279 14278 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14238 35199 14278 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 6042 14273 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5956 14273 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5870 14273 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5784 14273 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5698 14273 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5612 14273 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5526 14273 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5440 14273 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5354 14273 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5268 14273 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14233 5182 14273 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39931 14198 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39850 14198 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39769 14198 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39688 14198 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39607 14198 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39526 14198 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39445 14198 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39364 14198 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39283 14198 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39202 14198 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39121 14198 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 39040 14198 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38959 14198 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38879 14198 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38799 14198 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38719 14198 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38639 14198 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38559 14198 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38479 14198 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38399 14198 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38319 14198 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38239 14198 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38159 14198 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 38079 14198 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37999 14198 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37919 14198 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37839 14198 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37759 14198 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37679 14198 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37599 14198 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37519 14198 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37439 14198 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37359 14198 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37279 14198 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37199 14198 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37119 14198 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 37039 14198 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36959 14198 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36879 14198 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36799 14198 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36719 14198 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36639 14198 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36559 14198 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36479 14198 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36399 14198 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36319 14198 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36239 14198 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36159 14198 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 36079 14198 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35999 14198 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35919 14198 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35839 14198 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35759 14198 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35679 14198 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35599 14198 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35519 14198 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35439 14198 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35359 14198 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35279 14198 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14158 35199 14198 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 6042 14192 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5956 14192 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5870 14192 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5784 14192 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5698 14192 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5612 14192 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5526 14192 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5440 14192 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5354 14192 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5268 14192 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14152 5182 14192 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39931 14118 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39850 14118 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39769 14118 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39688 14118 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39607 14118 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39526 14118 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39445 14118 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39364 14118 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39283 14118 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39202 14118 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39121 14118 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 39040 14118 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38959 14118 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38879 14118 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38799 14118 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38719 14118 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38639 14118 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38559 14118 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38479 14118 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38399 14118 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38319 14118 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38239 14118 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38159 14118 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 38079 14118 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37999 14118 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37919 14118 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37839 14118 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37759 14118 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37679 14118 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37599 14118 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37519 14118 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37439 14118 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37359 14118 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37279 14118 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37199 14118 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37119 14118 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 37039 14118 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36959 14118 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36879 14118 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36799 14118 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36719 14118 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36639 14118 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36559 14118 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36479 14118 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36399 14118 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36319 14118 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36239 14118 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36159 14118 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 36079 14118 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35999 14118 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35919 14118 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35839 14118 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35759 14118 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35679 14118 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35599 14118 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35519 14118 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35439 14118 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35359 14118 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35279 14118 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14078 35199 14118 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 6042 14111 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5956 14111 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5870 14111 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5784 14111 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5698 14111 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5612 14111 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5526 14111 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5440 14111 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5354 14111 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5268 14111 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 14071 5182 14111 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39931 14038 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39850 14038 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39769 14038 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39688 14038 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39607 14038 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39526 14038 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39445 14038 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39364 14038 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39283 14038 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39202 14038 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39121 14038 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 39040 14038 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38959 14038 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38879 14038 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38799 14038 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38719 14038 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38639 14038 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38559 14038 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38479 14038 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38399 14038 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38319 14038 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38239 14038 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38159 14038 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 38079 14038 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37999 14038 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37919 14038 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37839 14038 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37759 14038 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37679 14038 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37599 14038 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37519 14038 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37439 14038 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37359 14038 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37279 14038 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37199 14038 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37119 14038 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 37039 14038 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36959 14038 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36879 14038 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36799 14038 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36719 14038 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36639 14038 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36559 14038 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36479 14038 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36399 14038 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36319 14038 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36239 14038 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36159 14038 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 36079 14038 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35999 14038 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35919 14038 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35839 14038 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35759 14038 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35679 14038 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35599 14038 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35519 14038 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35439 14038 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35359 14038 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35279 14038 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13998 35199 14038 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 6042 14030 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5956 14030 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5870 14030 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5784 14030 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5698 14030 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5612 14030 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5526 14030 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5440 14030 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5354 14030 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5268 14030 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13990 5182 14030 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39931 13958 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39850 13958 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39769 13958 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39688 13958 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39607 13958 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39526 13958 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39445 13958 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39364 13958 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39283 13958 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39202 13958 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39121 13958 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 39040 13958 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38959 13958 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38879 13958 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38799 13958 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38719 13958 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38639 13958 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38559 13958 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38479 13958 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38399 13958 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38319 13958 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38239 13958 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38159 13958 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 38079 13958 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37999 13958 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37919 13958 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37839 13958 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37759 13958 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37679 13958 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37599 13958 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37519 13958 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37439 13958 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37359 13958 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37279 13958 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37199 13958 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37119 13958 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 37039 13958 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36959 13958 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36879 13958 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36799 13958 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36719 13958 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36639 13958 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36559 13958 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36479 13958 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36399 13958 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36319 13958 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36239 13958 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36159 13958 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 36079 13958 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35999 13958 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35919 13958 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35839 13958 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35759 13958 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35679 13958 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35599 13958 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35519 13958 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35439 13958 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35359 13958 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35279 13958 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13918 35199 13958 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 6042 13949 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5956 13949 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5870 13949 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5784 13949 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5698 13949 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5612 13949 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5526 13949 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5440 13949 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5354 13949 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5268 13949 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13909 5182 13949 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39931 13878 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39850 13878 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39769 13878 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39688 13878 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39607 13878 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39526 13878 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39445 13878 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39364 13878 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39283 13878 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39202 13878 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39121 13878 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 39040 13878 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38959 13878 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38879 13878 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38799 13878 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38719 13878 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38639 13878 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38559 13878 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38479 13878 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38399 13878 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38319 13878 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38239 13878 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38159 13878 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 38079 13878 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37999 13878 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37919 13878 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37839 13878 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37759 13878 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37679 13878 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37599 13878 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37519 13878 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37439 13878 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37359 13878 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37279 13878 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37199 13878 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37119 13878 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 37039 13878 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36959 13878 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36879 13878 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36799 13878 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36719 13878 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36639 13878 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36559 13878 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36479 13878 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36399 13878 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36319 13878 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36239 13878 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36159 13878 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 36079 13878 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35999 13878 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35919 13878 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35839 13878 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35759 13878 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35679 13878 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35599 13878 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35519 13878 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35439 13878 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35359 13878 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35279 13878 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13838 35199 13878 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 6042 13868 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5956 13868 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5870 13868 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5784 13868 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5698 13868 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5612 13868 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5526 13868 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5440 13868 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5354 13868 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5268 13868 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13828 5182 13868 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39931 13798 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39850 13798 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39769 13798 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39688 13798 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39607 13798 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39526 13798 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39445 13798 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39364 13798 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39283 13798 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39202 13798 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39121 13798 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 39040 13798 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38959 13798 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38879 13798 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38799 13798 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38719 13798 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38639 13798 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38559 13798 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38479 13798 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38399 13798 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38319 13798 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38239 13798 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38159 13798 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 38079 13798 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37999 13798 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37919 13798 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37839 13798 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37759 13798 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37679 13798 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37599 13798 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37519 13798 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37439 13798 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37359 13798 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37279 13798 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37199 13798 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37119 13798 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 37039 13798 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36959 13798 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36879 13798 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36799 13798 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36719 13798 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36639 13798 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36559 13798 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36479 13798 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36399 13798 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36319 13798 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36239 13798 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36159 13798 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 36079 13798 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35999 13798 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35919 13798 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35839 13798 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35759 13798 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35679 13798 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35599 13798 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35519 13798 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35439 13798 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35359 13798 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35279 13798 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13758 35199 13798 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 6042 13787 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5956 13787 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5870 13787 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5784 13787 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5698 13787 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5612 13787 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5526 13787 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5440 13787 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5354 13787 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5268 13787 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13747 5182 13787 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39931 13718 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39850 13718 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39769 13718 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39688 13718 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39607 13718 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39526 13718 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39445 13718 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39364 13718 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39283 13718 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39202 13718 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39121 13718 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 39040 13718 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38959 13718 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38879 13718 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38799 13718 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38719 13718 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38639 13718 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38559 13718 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38479 13718 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38399 13718 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38319 13718 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38239 13718 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38159 13718 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 38079 13718 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37999 13718 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37919 13718 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37839 13718 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37759 13718 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37679 13718 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37599 13718 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37519 13718 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37439 13718 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37359 13718 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37279 13718 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37199 13718 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37119 13718 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 37039 13718 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36959 13718 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36879 13718 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36799 13718 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36719 13718 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36639 13718 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36559 13718 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36479 13718 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36399 13718 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36319 13718 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36239 13718 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36159 13718 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 36079 13718 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35999 13718 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35919 13718 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35839 13718 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35759 13718 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35679 13718 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35599 13718 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35519 13718 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35439 13718 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35359 13718 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35279 13718 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13678 35199 13718 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 6042 13706 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5956 13706 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5870 13706 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5784 13706 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5698 13706 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5612 13706 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5526 13706 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5440 13706 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5354 13706 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5268 13706 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13666 5182 13706 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39931 13638 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39850 13638 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39769 13638 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39688 13638 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39607 13638 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39526 13638 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39445 13638 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39364 13638 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39283 13638 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39202 13638 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39121 13638 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 39040 13638 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38959 13638 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38879 13638 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38799 13638 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38719 13638 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38639 13638 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38559 13638 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38479 13638 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38399 13638 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38319 13638 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38239 13638 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38159 13638 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 38079 13638 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37999 13638 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37919 13638 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37839 13638 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37759 13638 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37679 13638 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37599 13638 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37519 13638 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37439 13638 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37359 13638 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37279 13638 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37199 13638 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37119 13638 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 37039 13638 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36959 13638 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36879 13638 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36799 13638 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36719 13638 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36639 13638 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36559 13638 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36479 13638 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36399 13638 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36319 13638 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36239 13638 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36159 13638 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 36079 13638 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35999 13638 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35919 13638 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35839 13638 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35759 13638 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35679 13638 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35599 13638 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35519 13638 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35439 13638 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35359 13638 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35279 13638 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13598 35199 13638 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 6042 13625 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5956 13625 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5870 13625 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5784 13625 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5698 13625 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5612 13625 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5526 13625 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5440 13625 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5354 13625 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5268 13625 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13585 5182 13625 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39931 13558 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39850 13558 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39769 13558 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39688 13558 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39607 13558 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39526 13558 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39445 13558 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39364 13558 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39283 13558 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39202 13558 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39121 13558 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 39040 13558 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38959 13558 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38879 13558 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38799 13558 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38719 13558 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38639 13558 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38559 13558 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38479 13558 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38399 13558 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38319 13558 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38239 13558 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38159 13558 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 38079 13558 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37999 13558 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37919 13558 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37839 13558 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37759 13558 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37679 13558 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37599 13558 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37519 13558 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37439 13558 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37359 13558 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37279 13558 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37199 13558 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37119 13558 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 37039 13558 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36959 13558 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36879 13558 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36799 13558 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36719 13558 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36639 13558 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36559 13558 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36479 13558 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36399 13558 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36319 13558 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36239 13558 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36159 13558 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 36079 13558 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35999 13558 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35919 13558 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35839 13558 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35759 13558 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35679 13558 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35599 13558 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35519 13558 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35439 13558 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35359 13558 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35279 13558 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13518 35199 13558 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 6042 13544 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5956 13544 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5870 13544 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5784 13544 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5698 13544 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5612 13544 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5526 13544 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5440 13544 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5354 13544 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5268 13544 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13504 5182 13544 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39931 13478 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39850 13478 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39769 13478 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39688 13478 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39607 13478 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39526 13478 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39445 13478 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39364 13478 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39283 13478 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39202 13478 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39121 13478 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 39040 13478 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38959 13478 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38879 13478 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38799 13478 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38719 13478 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38639 13478 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38559 13478 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38479 13478 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38399 13478 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38319 13478 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38239 13478 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38159 13478 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 38079 13478 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37999 13478 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37919 13478 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37839 13478 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37759 13478 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37679 13478 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37599 13478 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37519 13478 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37439 13478 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37359 13478 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37279 13478 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37199 13478 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37119 13478 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 37039 13478 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36959 13478 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36879 13478 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36799 13478 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36719 13478 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36639 13478 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36559 13478 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36479 13478 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36399 13478 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36319 13478 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36239 13478 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36159 13478 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 36079 13478 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35999 13478 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35919 13478 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35839 13478 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35759 13478 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35679 13478 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35599 13478 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35519 13478 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35439 13478 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35359 13478 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35279 13478 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13438 35199 13478 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 6042 13463 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5956 13463 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5870 13463 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5784 13463 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5698 13463 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5612 13463 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5526 13463 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5440 13463 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5354 13463 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5268 13463 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13423 5182 13463 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39931 13398 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39850 13398 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39769 13398 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39688 13398 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39607 13398 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39526 13398 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39445 13398 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39364 13398 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39283 13398 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39202 13398 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39121 13398 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 39040 13398 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38959 13398 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38879 13398 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38799 13398 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38719 13398 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38639 13398 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38559 13398 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38479 13398 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38399 13398 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38319 13398 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38239 13398 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38159 13398 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 38079 13398 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37999 13398 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37919 13398 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37839 13398 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37759 13398 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37679 13398 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37599 13398 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37519 13398 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37439 13398 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37359 13398 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37279 13398 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37199 13398 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37119 13398 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 37039 13398 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36959 13398 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36879 13398 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36799 13398 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36719 13398 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36639 13398 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36559 13398 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36479 13398 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36399 13398 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36319 13398 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36239 13398 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36159 13398 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 36079 13398 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35999 13398 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35919 13398 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35839 13398 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35759 13398 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35679 13398 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35599 13398 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35519 13398 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35439 13398 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35359 13398 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35279 13398 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13358 35199 13398 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 6042 13382 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5956 13382 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5870 13382 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5784 13382 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5698 13382 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5612 13382 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5526 13382 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5440 13382 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5354 13382 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5268 13382 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13342 5182 13382 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39931 13318 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39850 13318 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39769 13318 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39688 13318 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39607 13318 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39526 13318 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39445 13318 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39364 13318 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39283 13318 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39202 13318 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39121 13318 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 39040 13318 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38959 13318 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38879 13318 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38799 13318 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38719 13318 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38639 13318 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38559 13318 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38479 13318 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38399 13318 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38319 13318 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38239 13318 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38159 13318 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 38079 13318 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37999 13318 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37919 13318 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37839 13318 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37759 13318 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37679 13318 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37599 13318 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37519 13318 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37439 13318 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37359 13318 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37279 13318 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37199 13318 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37119 13318 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 37039 13318 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36959 13318 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36879 13318 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36799 13318 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36719 13318 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36639 13318 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36559 13318 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36479 13318 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36399 13318 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36319 13318 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36239 13318 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36159 13318 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 36079 13318 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35999 13318 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35919 13318 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35839 13318 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35759 13318 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35679 13318 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35599 13318 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35519 13318 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35439 13318 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35359 13318 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35279 13318 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13278 35199 13318 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 6042 13301 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5956 13301 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5870 13301 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5784 13301 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5698 13301 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5612 13301 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5526 13301 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5440 13301 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5354 13301 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5268 13301 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13261 5182 13301 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39931 13238 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39850 13238 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39769 13238 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39688 13238 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39607 13238 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39526 13238 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39445 13238 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39364 13238 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39283 13238 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39202 13238 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39121 13238 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 39040 13238 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38959 13238 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38879 13238 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38799 13238 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38719 13238 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38639 13238 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38559 13238 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38479 13238 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38399 13238 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38319 13238 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38239 13238 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38159 13238 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 38079 13238 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37999 13238 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37919 13238 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37839 13238 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37759 13238 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37679 13238 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37599 13238 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37519 13238 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37439 13238 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37359 13238 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37279 13238 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37199 13238 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37119 13238 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 37039 13238 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36959 13238 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36879 13238 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36799 13238 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36719 13238 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36639 13238 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36559 13238 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36479 13238 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36399 13238 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36319 13238 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36239 13238 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36159 13238 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 36079 13238 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35999 13238 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35919 13238 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35839 13238 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35759 13238 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35679 13238 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35599 13238 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35519 13238 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35439 13238 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35359 13238 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35279 13238 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13198 35199 13238 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 6042 13220 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5956 13220 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5870 13220 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5784 13220 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5698 13220 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5612 13220 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5526 13220 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5440 13220 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5354 13220 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5268 13220 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13180 5182 13220 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39931 13158 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39850 13158 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39769 13158 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39688 13158 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39607 13158 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39526 13158 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39445 13158 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39364 13158 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39283 13158 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39202 13158 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39121 13158 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 39040 13158 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38959 13158 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38879 13158 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38799 13158 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38719 13158 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38639 13158 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38559 13158 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38479 13158 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38399 13158 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38319 13158 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38239 13158 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38159 13158 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 38079 13158 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37999 13158 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37919 13158 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37839 13158 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37759 13158 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37679 13158 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37599 13158 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37519 13158 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37439 13158 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37359 13158 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37279 13158 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37199 13158 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37119 13158 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 37039 13158 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36959 13158 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36879 13158 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36799 13158 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36719 13158 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36639 13158 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36559 13158 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36479 13158 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36399 13158 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36319 13158 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36239 13158 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36159 13158 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 36079 13158 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35999 13158 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35919 13158 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35839 13158 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35759 13158 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35679 13158 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35599 13158 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35519 13158 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35439 13158 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35359 13158 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35279 13158 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13118 35199 13158 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 6042 13139 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5956 13139 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5870 13139 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5784 13139 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5698 13139 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5612 13139 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5526 13139 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5440 13139 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5354 13139 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5268 13139 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13099 5182 13139 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39931 13078 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39850 13078 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39769 13078 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39688 13078 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39607 13078 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39526 13078 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39445 13078 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39364 13078 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39283 13078 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39202 13078 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39121 13078 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 39040 13078 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38959 13078 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38879 13078 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38799 13078 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38719 13078 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38639 13078 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38559 13078 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38479 13078 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38399 13078 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38319 13078 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38239 13078 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38159 13078 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 38079 13078 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37999 13078 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37919 13078 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37839 13078 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37759 13078 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37679 13078 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37599 13078 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37519 13078 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37439 13078 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37359 13078 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37279 13078 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37199 13078 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37119 13078 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 37039 13078 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36959 13078 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36879 13078 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36799 13078 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36719 13078 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36639 13078 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36559 13078 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36479 13078 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36399 13078 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36319 13078 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36239 13078 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36159 13078 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 36079 13078 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35999 13078 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35919 13078 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35839 13078 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35759 13078 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35679 13078 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35599 13078 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35519 13078 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35439 13078 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35359 13078 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35279 13078 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13038 35199 13078 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 6042 13058 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5956 13058 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5870 13058 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5784 13058 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5698 13058 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5612 13058 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5526 13058 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5440 13058 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5354 13058 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5268 13058 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 13018 5182 13058 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39931 12998 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39850 12998 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39769 12998 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39688 12998 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39607 12998 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39526 12998 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39445 12998 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39364 12998 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39283 12998 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39202 12998 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39121 12998 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 39040 12998 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38959 12998 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38879 12998 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38799 12998 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38719 12998 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38639 12998 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38559 12998 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38479 12998 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38399 12998 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38319 12998 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38239 12998 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38159 12998 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 38079 12998 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37999 12998 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37919 12998 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37839 12998 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37759 12998 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37679 12998 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37599 12998 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37519 12998 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37439 12998 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37359 12998 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37279 12998 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37199 12998 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37119 12998 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 37039 12998 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36959 12998 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36879 12998 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36799 12998 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36719 12998 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36639 12998 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36559 12998 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36479 12998 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36399 12998 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36319 12998 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36239 12998 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36159 12998 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 36079 12998 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35999 12998 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35919 12998 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35839 12998 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35759 12998 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35679 12998 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35599 12998 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35519 12998 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35439 12998 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35359 12998 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35279 12998 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12958 35199 12998 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 6042 12977 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5956 12977 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5870 12977 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5784 12977 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5698 12977 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5612 12977 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5526 12977 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5440 12977 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5354 12977 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5268 12977 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12937 5182 12977 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39931 12918 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39850 12918 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39769 12918 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39688 12918 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39607 12918 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39526 12918 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39445 12918 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39364 12918 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39283 12918 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39202 12918 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39121 12918 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 39040 12918 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38959 12918 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38879 12918 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38799 12918 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38719 12918 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38639 12918 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38559 12918 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38479 12918 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38399 12918 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38319 12918 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38239 12918 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38159 12918 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 38079 12918 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37999 12918 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37919 12918 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37839 12918 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37759 12918 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37679 12918 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37599 12918 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37519 12918 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37439 12918 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37359 12918 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37279 12918 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37199 12918 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37119 12918 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 37039 12918 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36959 12918 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36879 12918 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36799 12918 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36719 12918 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36639 12918 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36559 12918 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36479 12918 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36399 12918 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36319 12918 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36239 12918 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36159 12918 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 36079 12918 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35999 12918 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35919 12918 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35839 12918 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35759 12918 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35679 12918 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35599 12918 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35519 12918 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35439 12918 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35359 12918 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35279 12918 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12878 35199 12918 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 6042 12896 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5956 12896 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5870 12896 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5784 12896 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5698 12896 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5612 12896 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5526 12896 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5440 12896 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5354 12896 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5268 12896 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12856 5182 12896 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39931 12838 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39850 12838 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39769 12838 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39688 12838 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39607 12838 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39526 12838 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39445 12838 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39364 12838 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39283 12838 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39202 12838 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39121 12838 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 39040 12838 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38959 12838 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38879 12838 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38799 12838 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38719 12838 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38639 12838 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38559 12838 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38479 12838 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38399 12838 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38319 12838 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38239 12838 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38159 12838 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 38079 12838 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37999 12838 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37919 12838 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37839 12838 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37759 12838 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37679 12838 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37599 12838 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37519 12838 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37439 12838 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37359 12838 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37279 12838 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37199 12838 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37119 12838 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 37039 12838 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36959 12838 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36879 12838 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36799 12838 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36719 12838 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36639 12838 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36559 12838 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36479 12838 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36399 12838 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36319 12838 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36239 12838 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36159 12838 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 36079 12838 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35999 12838 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35919 12838 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35839 12838 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35759 12838 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35679 12838 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35599 12838 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35519 12838 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35439 12838 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35359 12838 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35279 12838 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12798 35199 12838 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 6042 12815 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5956 12815 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5870 12815 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5784 12815 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5698 12815 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5612 12815 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5526 12815 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5440 12815 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5354 12815 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5268 12815 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12775 5182 12815 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39931 12758 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39850 12758 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39769 12758 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39688 12758 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39607 12758 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39526 12758 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39445 12758 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39364 12758 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39283 12758 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39202 12758 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39121 12758 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 39040 12758 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38959 12758 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38879 12758 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38799 12758 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38719 12758 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38639 12758 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38559 12758 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38479 12758 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38399 12758 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38319 12758 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38239 12758 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38159 12758 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 38079 12758 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37999 12758 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37919 12758 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37839 12758 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37759 12758 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37679 12758 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37599 12758 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37519 12758 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37439 12758 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37359 12758 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37279 12758 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37199 12758 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37119 12758 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 37039 12758 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36959 12758 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36879 12758 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36799 12758 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36719 12758 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36639 12758 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36559 12758 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36479 12758 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36399 12758 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36319 12758 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36239 12758 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36159 12758 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 36079 12758 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35999 12758 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35919 12758 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35839 12758 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35759 12758 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35679 12758 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35599 12758 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35519 12758 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35439 12758 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35359 12758 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35279 12758 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12718 35199 12758 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 6042 12734 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5956 12734 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5870 12734 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5784 12734 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5698 12734 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5612 12734 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5526 12734 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5440 12734 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5354 12734 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5268 12734 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12694 5182 12734 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39931 12678 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39850 12678 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39769 12678 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39688 12678 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39607 12678 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39526 12678 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39445 12678 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39364 12678 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39283 12678 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39202 12678 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39121 12678 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 39040 12678 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38959 12678 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38879 12678 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38799 12678 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38719 12678 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38639 12678 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38559 12678 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38479 12678 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38399 12678 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38319 12678 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38239 12678 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38159 12678 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 38079 12678 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37999 12678 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37919 12678 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37839 12678 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37759 12678 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37679 12678 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37599 12678 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37519 12678 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37439 12678 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37359 12678 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37279 12678 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37199 12678 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37119 12678 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 37039 12678 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36959 12678 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36879 12678 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36799 12678 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36719 12678 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36639 12678 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36559 12678 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36479 12678 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36399 12678 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36319 12678 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36239 12678 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36159 12678 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 36079 12678 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35999 12678 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35919 12678 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35839 12678 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35759 12678 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35679 12678 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35599 12678 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35519 12678 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35439 12678 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35359 12678 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35279 12678 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12638 35199 12678 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 6042 12653 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5956 12653 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5870 12653 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5784 12653 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5698 12653 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5612 12653 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5526 12653 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5440 12653 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5354 12653 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5268 12653 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12613 5182 12653 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39931 12598 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39850 12598 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39769 12598 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39688 12598 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39607 12598 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39526 12598 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39445 12598 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39364 12598 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39283 12598 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39202 12598 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39121 12598 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 39040 12598 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38959 12598 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38879 12598 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38799 12598 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38719 12598 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38639 12598 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38559 12598 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38479 12598 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38399 12598 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38319 12598 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38239 12598 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38159 12598 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 38079 12598 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37999 12598 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37919 12598 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37839 12598 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37759 12598 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37679 12598 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37599 12598 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37519 12598 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37439 12598 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37359 12598 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37279 12598 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37199 12598 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37119 12598 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 37039 12598 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36959 12598 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36879 12598 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36799 12598 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36719 12598 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36639 12598 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36559 12598 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36479 12598 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36399 12598 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36319 12598 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36239 12598 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36159 12598 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 36079 12598 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35999 12598 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35919 12598 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35839 12598 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35759 12598 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35679 12598 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35599 12598 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35519 12598 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35439 12598 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35359 12598 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35279 12598 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12558 35199 12598 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 6042 12572 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5956 12572 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5870 12572 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5784 12572 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5698 12572 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5612 12572 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5526 12572 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5440 12572 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5354 12572 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5268 12572 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12532 5182 12572 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39931 12518 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39850 12518 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39769 12518 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39688 12518 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39607 12518 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39526 12518 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39445 12518 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39364 12518 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39283 12518 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39202 12518 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39121 12518 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 39040 12518 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38959 12518 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38879 12518 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38799 12518 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38719 12518 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38639 12518 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38559 12518 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38479 12518 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38399 12518 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38319 12518 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38239 12518 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38159 12518 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 38079 12518 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37999 12518 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37919 12518 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37839 12518 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37759 12518 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37679 12518 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37599 12518 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37519 12518 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37439 12518 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37359 12518 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37279 12518 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37199 12518 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37119 12518 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 37039 12518 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36959 12518 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36879 12518 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36799 12518 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36719 12518 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36639 12518 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36559 12518 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36479 12518 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36399 12518 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36319 12518 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36239 12518 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36159 12518 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 36079 12518 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35999 12518 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35919 12518 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35839 12518 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35759 12518 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35679 12518 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35599 12518 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35519 12518 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35439 12518 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35359 12518 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35279 12518 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12478 35199 12518 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 6042 12491 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5956 12491 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5870 12491 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5784 12491 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5698 12491 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5612 12491 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5526 12491 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5440 12491 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5354 12491 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5268 12491 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12451 5182 12491 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39931 12438 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39850 12438 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39769 12438 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39688 12438 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39607 12438 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39526 12438 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39445 12438 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39364 12438 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39283 12438 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39202 12438 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39121 12438 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 39040 12438 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38959 12438 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38879 12438 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38799 12438 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38719 12438 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38639 12438 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38559 12438 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38479 12438 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38399 12438 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38319 12438 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38239 12438 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38159 12438 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 38079 12438 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37999 12438 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37919 12438 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37839 12438 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37759 12438 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37679 12438 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37599 12438 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37519 12438 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37439 12438 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37359 12438 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37279 12438 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37199 12438 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37119 12438 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 37039 12438 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36959 12438 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36879 12438 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36799 12438 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36719 12438 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36639 12438 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36559 12438 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36479 12438 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36399 12438 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36319 12438 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36239 12438 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36159 12438 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 36079 12438 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35999 12438 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35919 12438 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35839 12438 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35759 12438 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35679 12438 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35599 12438 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35519 12438 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35439 12438 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35359 12438 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35279 12438 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12398 35199 12438 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 6042 12410 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5956 12410 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5870 12410 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5784 12410 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5698 12410 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5612 12410 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5526 12410 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5440 12410 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5354 12410 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5268 12410 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12370 5182 12410 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39931 12358 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39850 12358 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39769 12358 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39688 12358 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39607 12358 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39526 12358 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39445 12358 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39364 12358 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39283 12358 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39202 12358 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39121 12358 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 39040 12358 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38959 12358 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38879 12358 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38799 12358 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38719 12358 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38639 12358 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38559 12358 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38479 12358 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38399 12358 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38319 12358 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38239 12358 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38159 12358 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 38079 12358 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37999 12358 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37919 12358 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37839 12358 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37759 12358 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37679 12358 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37599 12358 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37519 12358 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37439 12358 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37359 12358 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37279 12358 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37199 12358 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37119 12358 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 37039 12358 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36959 12358 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36879 12358 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36799 12358 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36719 12358 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36639 12358 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36559 12358 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36479 12358 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36399 12358 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36319 12358 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36239 12358 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36159 12358 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 36079 12358 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35999 12358 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35919 12358 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35839 12358 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35759 12358 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35679 12358 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35599 12358 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35519 12358 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35439 12358 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35359 12358 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35279 12358 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12318 35199 12358 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 6042 12329 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5956 12329 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5870 12329 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5784 12329 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5698 12329 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5612 12329 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5526 12329 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5440 12329 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5354 12329 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5268 12329 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12289 5182 12329 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12212 39930 12252 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12212 39850 12252 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12212 39770 12252 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12212 39690 12252 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12212 39610 12252 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12212 39530 12252 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12212 39450 12252 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 6042 12248 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5956 12248 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5870 12248 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5784 12248 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5698 12248 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5612 12248 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5526 12248 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5440 12248 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5354 12248 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5268 12248 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12208 5182 12248 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12182 39341 12222 39381 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12182 39259 12222 39299 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12132 39930 12172 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12132 39850 12172 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12132 39770 12172 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12132 39690 12172 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12132 39610 12172 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12132 39530 12172 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12132 39450 12172 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 6042 12167 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5956 12167 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5870 12167 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5784 12167 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5698 12167 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5612 12167 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5526 12167 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5440 12167 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5354 12167 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5268 12167 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12127 5182 12167 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12052 39930 12092 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12052 39850 12092 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12052 39770 12092 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12052 39690 12092 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12052 39610 12092 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12052 39530 12092 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12052 39450 12092 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 6042 12086 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5956 12086 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5870 12086 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5784 12086 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5698 12086 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5612 12086 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5526 12086 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5440 12086 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5354 12086 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5268 12086 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 12046 5182 12086 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11972 39930 12012 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11972 39850 12012 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11972 39770 12012 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11972 39690 12012 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11972 39610 12012 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11972 39530 12012 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11972 39450 12012 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 6042 12005 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5956 12005 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5870 12005 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5784 12005 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5698 12005 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5612 12005 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5526 12005 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5440 12005 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5354 12005 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5268 12005 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11965 5182 12005 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11892 39930 11932 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11892 39850 11932 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11892 39770 11932 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11892 39690 11932 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11892 39610 11932 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11892 39530 11932 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11892 39450 11932 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 6042 11924 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5956 11924 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5870 11924 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5784 11924 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5698 11924 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5612 11924 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5526 11924 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5440 11924 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5354 11924 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5268 11924 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11884 5182 11924 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11812 39930 11852 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11812 39850 11852 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11812 39770 11852 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11812 39690 11852 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11812 39610 11852 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11812 39530 11852 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11812 39450 11852 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 6042 11843 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5956 11843 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5870 11843 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5784 11843 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5698 11843 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5612 11843 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5526 11843 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5440 11843 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5354 11843 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5268 11843 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11803 5182 11843 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11732 39930 11772 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11732 39850 11772 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11732 39770 11772 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11732 39690 11772 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11732 39610 11772 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11732 39530 11772 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11732 39450 11772 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 6042 11762 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5956 11762 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5870 11762 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5784 11762 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5698 11762 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5612 11762 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5526 11762 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5440 11762 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5354 11762 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5268 11762 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11722 5182 11762 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11652 39930 11692 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11652 39850 11692 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11652 39770 11692 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11652 39690 11692 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11652 39610 11692 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11652 39530 11692 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11652 39450 11692 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 6042 11681 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5956 11681 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5870 11681 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5784 11681 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5698 11681 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5612 11681 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5526 11681 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5440 11681 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5354 11681 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5268 11681 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11641 5182 11681 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11572 39930 11612 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11572 39850 11612 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11572 39770 11612 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11572 39690 11612 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11572 39610 11612 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11572 39530 11612 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11572 39450 11612 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 6042 11600 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5956 11600 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5870 11600 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5784 11600 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5698 11600 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5612 11600 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5526 11600 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5440 11600 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5354 11600 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5268 11600 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11560 5182 11600 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11492 39930 11532 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11492 39850 11532 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11492 39770 11532 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11492 39690 11532 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11492 39610 11532 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11492 39530 11532 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11492 39450 11532 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 6042 11519 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5956 11519 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5870 11519 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5784 11519 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5698 11519 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5612 11519 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5526 11519 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5440 11519 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5354 11519 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5268 11519 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11479 5182 11519 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11412 39930 11452 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11412 39850 11452 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11412 39770 11452 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11412 39690 11452 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11412 39610 11452 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11412 39530 11452 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11412 39450 11452 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 6042 11438 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5956 11438 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5870 11438 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5784 11438 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5698 11438 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5612 11438 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5526 11438 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5440 11438 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5354 11438 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5268 11438 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11398 5182 11438 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11332 39930 11372 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11332 39850 11372 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11332 39770 11372 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11332 39690 11372 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11332 39610 11372 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11332 39530 11372 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11332 39450 11372 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 6042 11357 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5956 11357 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5870 11357 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5784 11357 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5698 11357 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5612 11357 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5526 11357 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5440 11357 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5354 11357 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5268 11357 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11317 5182 11357 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11252 39930 11292 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11252 39850 11292 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11252 39770 11292 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11252 39690 11292 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11252 39610 11292 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11252 39530 11292 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11252 39450 11292 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 6042 11276 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5956 11276 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5870 11276 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5784 11276 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5698 11276 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5612 11276 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5526 11276 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5440 11276 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5354 11276 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5268 11276 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11236 5182 11276 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11172 39930 11212 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11172 39850 11212 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11172 39770 11212 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11172 39690 11212 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11172 39610 11212 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11172 39530 11212 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11172 39450 11212 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 6042 11195 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5956 11195 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5870 11195 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5784 11195 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5698 11195 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5612 11195 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5526 11195 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5440 11195 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5354 11195 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5268 11195 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11155 5182 11195 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11092 39930 11132 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11092 39850 11132 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11092 39770 11132 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11092 39690 11132 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11092 39610 11132 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11092 39530 11132 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11092 39450 11132 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 6042 11114 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5956 11114 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5870 11114 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5784 11114 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5698 11114 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5612 11114 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5526 11114 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5440 11114 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5354 11114 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5268 11114 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11074 5182 11114 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11012 39930 11052 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11012 39850 11052 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11012 39770 11052 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11012 39690 11052 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11012 39610 11052 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11012 39530 11052 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 11012 39450 11052 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 6042 11033 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5956 11033 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5870 11033 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5784 11033 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5698 11033 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5612 11033 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5526 11033 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5440 11033 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5354 11033 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5268 11033 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10993 5182 11033 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10932 39930 10972 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10932 39850 10972 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10932 39770 10972 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10932 39690 10972 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10932 39610 10972 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10932 39530 10972 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10932 39450 10972 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 6042 10952 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5956 10952 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5870 10952 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5784 10952 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5698 10952 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5612 10952 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5526 10952 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5440 10952 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5354 10952 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5268 10952 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10912 5182 10952 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10852 39930 10892 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10852 39850 10892 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10852 39770 10892 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10852 39690 10892 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10852 39610 10892 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10852 39530 10892 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10852 39450 10892 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 6042 10871 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5956 10871 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5870 10871 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5784 10871 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5698 10871 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5612 10871 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5526 10871 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5440 10871 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5354 10871 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5268 10871 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10831 5182 10871 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10772 39930 10812 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10772 39850 10812 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10772 39770 10812 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10772 39690 10812 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10772 39610 10812 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10772 39530 10812 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10772 39450 10812 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 6042 10790 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5956 10790 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5870 10790 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5784 10790 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5698 10790 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5612 10790 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5526 10790 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5440 10790 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5354 10790 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5268 10790 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10750 5182 10790 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10692 39930 10732 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10692 39850 10732 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10692 39770 10732 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10692 39690 10732 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10692 39610 10732 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10692 39530 10732 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10692 39450 10732 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 6042 10709 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5956 10709 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5870 10709 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5784 10709 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5698 10709 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5612 10709 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5526 10709 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5440 10709 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5354 10709 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5268 10709 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10669 5182 10709 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10612 39930 10652 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10612 39850 10652 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10612 39770 10652 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10612 39690 10652 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10612 39610 10652 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10612 39530 10652 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10612 39450 10652 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 6042 10628 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5956 10628 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5870 10628 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5784 10628 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5698 10628 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5612 10628 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5526 10628 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5440 10628 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5354 10628 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5268 10628 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10588 5182 10628 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10532 39930 10572 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10532 39850 10572 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10532 39770 10572 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10532 39690 10572 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10532 39610 10572 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10532 39530 10572 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10532 39450 10572 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 6042 10546 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5956 10546 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5870 10546 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5784 10546 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5698 10546 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5612 10546 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5526 10546 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5440 10546 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5354 10546 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5268 10546 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10506 5182 10546 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10452 39930 10492 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10452 39850 10492 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10452 39770 10492 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10452 39690 10492 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10452 39610 10492 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10452 39530 10492 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10452 39450 10492 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 6042 10464 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5956 10464 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5870 10464 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5784 10464 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5698 10464 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5612 10464 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5526 10464 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5440 10464 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5354 10464 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5268 10464 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10424 5182 10464 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10372 39930 10412 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10372 39850 10412 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10372 39770 10412 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10372 39690 10412 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10372 39610 10412 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10372 39530 10412 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10372 39450 10412 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 6042 10382 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5956 10382 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5870 10382 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5784 10382 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5698 10382 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5612 10382 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5526 10382 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5440 10382 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5354 10382 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5268 10382 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10342 5182 10382 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10292 39930 10332 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10292 39850 10332 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10292 39770 10332 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10292 39690 10332 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10292 39610 10332 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10292 39530 10332 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10292 39450 10332 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 6042 10300 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5956 10300 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5870 10300 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5784 10300 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5698 10300 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5612 10300 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5526 10300 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5440 10300 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5354 10300 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5268 10300 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10260 5182 10300 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10212 39930 10252 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10212 39850 10252 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10212 39770 10252 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10212 39690 10252 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10212 39610 10252 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10212 39530 10252 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10212 39450 10252 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 6042 10218 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5956 10218 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5870 10218 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5784 10218 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5698 10218 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5612 10218 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5526 10218 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5440 10218 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5354 10218 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5268 10218 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10178 5182 10218 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10132 39930 10172 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10132 39850 10172 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10132 39770 10172 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10132 39690 10172 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10132 39610 10172 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10132 39530 10172 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10132 39450 10172 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 6042 10136 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5956 10136 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5870 10136 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5784 10136 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5698 10136 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5612 10136 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5526 10136 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5440 10136 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5354 10136 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5268 10136 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10096 5182 10136 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10052 39930 10092 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10052 39850 10092 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10052 39770 10092 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10052 39690 10092 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10052 39610 10092 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10052 39530 10092 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 10052 39450 10092 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9972 39930 10012 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9972 39850 10012 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9972 39770 10012 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9972 39690 10012 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9972 39610 10012 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9972 39530 10012 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9972 39450 10012 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9892 39930 9932 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9892 39850 9932 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9892 39770 9932 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9892 39690 9932 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9892 39610 9932 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9892 39530 9932 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9892 39450 9932 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9812 39930 9852 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9812 39850 9852 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9812 39770 9852 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9812 39690 9852 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9812 39610 9852 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9812 39530 9852 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9812 39450 9852 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9732 39930 9772 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9732 39850 9772 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9732 39770 9772 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9732 39690 9772 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9732 39610 9772 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9732 39530 9772 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9732 39450 9772 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9652 39930 9692 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9652 39850 9692 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9652 39770 9692 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9652 39690 9692 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9652 39610 9692 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9652 39530 9692 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9652 39450 9692 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9572 39930 9612 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9572 39850 9612 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9572 39770 9612 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9572 39690 9612 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9572 39610 9612 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9572 39530 9612 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9572 39450 9612 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9492 39930 9532 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9492 39850 9532 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9492 39770 9532 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9492 39690 9532 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9492 39610 9532 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9492 39530 9532 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9492 39450 9532 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9412 39930 9452 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9412 39850 9452 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9412 39770 9452 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9412 39690 9452 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9412 39610 9452 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9412 39530 9452 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9412 39450 9452 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9332 39930 9372 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9332 39850 9372 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9332 39770 9372 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9332 39690 9372 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9332 39610 9372 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9332 39530 9372 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9332 39450 9372 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9252 39930 9292 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9252 39850 9292 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9252 39770 9292 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9252 39690 9292 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9252 39610 9292 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9252 39530 9292 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9252 39450 9292 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9172 39930 9212 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9172 39850 9212 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9172 39770 9212 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9172 39690 9212 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9172 39610 9212 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9172 39530 9212 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9172 39450 9212 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9092 39930 9132 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9092 39850 9132 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9092 39770 9132 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9092 39690 9132 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9092 39610 9132 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9092 39530 9132 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9092 39450 9132 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9012 39930 9052 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9012 39850 9052 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9012 39770 9052 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9012 39690 9052 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9012 39610 9052 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9012 39530 9052 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 9012 39450 9052 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8932 39930 8972 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8932 39850 8972 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8932 39770 8972 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8932 39690 8972 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8932 39610 8972 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8932 39530 8972 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8932 39450 8972 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8852 39930 8892 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8852 39850 8892 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8852 39770 8892 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8852 39690 8892 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8852 39610 8892 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8852 39530 8892 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8852 39450 8892 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8772 39930 8812 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8772 39850 8812 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8772 39770 8812 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8772 39690 8812 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8772 39610 8812 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8772 39530 8812 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8772 39450 8812 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8692 39930 8732 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8692 39850 8732 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8692 39770 8732 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8692 39690 8732 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8692 39610 8732 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8692 39530 8732 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8692 39450 8732 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8612 39930 8652 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8612 39850 8652 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8612 39770 8652 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8612 39690 8652 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8612 39610 8652 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8612 39530 8652 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8612 39450 8652 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8532 39930 8572 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8532 39850 8572 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8532 39770 8572 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8532 39690 8572 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8532 39610 8572 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8532 39530 8572 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8532 39450 8572 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8452 39930 8492 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8452 39850 8492 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8452 39770 8492 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8452 39690 8492 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8452 39610 8492 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8452 39530 8492 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8452 39450 8492 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8372 39930 8412 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8372 39850 8412 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8372 39770 8412 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8372 39690 8412 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8372 39610 8412 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8372 39530 8412 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8372 39450 8412 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8292 39930 8332 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8292 39850 8332 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8292 39770 8332 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8292 39690 8332 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8292 39610 8332 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8292 39530 8332 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8292 39450 8332 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8212 39930 8252 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8212 39850 8252 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8212 39770 8252 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8212 39690 8252 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8212 39610 8252 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8212 39530 8252 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8212 39450 8252 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8132 39930 8172 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8132 39850 8172 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8132 39770 8172 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8132 39690 8172 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8132 39610 8172 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8132 39530 8172 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8132 39450 8172 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8052 39930 8092 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8052 39850 8092 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8052 39770 8092 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8052 39690 8092 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8052 39610 8092 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8052 39530 8092 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 8052 39450 8092 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7972 39930 8012 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7972 39850 8012 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7972 39770 8012 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7972 39690 8012 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7972 39610 8012 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7972 39530 8012 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7972 39450 8012 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7892 39930 7932 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7892 39850 7932 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7892 39770 7932 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7892 39690 7932 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7892 39610 7932 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7892 39530 7932 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7892 39450 7932 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7812 39930 7852 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7812 39850 7852 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7812 39770 7852 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7812 39690 7852 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7812 39610 7852 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7812 39530 7852 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7812 39450 7852 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7732 39930 7772 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7732 39850 7772 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7732 39770 7772 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7732 39690 7772 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7732 39610 7772 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7732 39530 7772 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7732 39450 7772 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7652 39930 7692 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7652 39850 7692 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7652 39770 7692 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7652 39690 7692 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7652 39610 7692 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7652 39530 7692 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7652 39450 7692 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7572 39930 7612 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7572 39850 7612 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7572 39770 7612 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7572 39690 7612 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7572 39610 7612 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7572 39530 7612 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7572 39450 7612 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7492 39930 7532 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7492 39850 7532 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7492 39770 7532 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7492 39690 7532 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7492 39610 7532 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7492 39530 7532 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7492 39450 7532 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7412 39930 7452 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7412 39850 7452 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7412 39770 7452 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7412 39690 7452 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7412 39610 7452 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7412 39530 7452 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7412 39450 7452 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7332 39930 7372 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7332 39850 7372 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7332 39770 7372 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7332 39690 7372 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7332 39610 7372 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7332 39530 7372 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7332 39450 7372 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7252 39930 7292 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7252 39850 7292 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7252 39770 7292 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7252 39690 7292 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7252 39610 7292 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7252 39530 7292 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7252 39450 7292 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7172 39930 7212 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7172 39850 7212 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7172 39770 7212 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7172 39690 7212 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7172 39610 7212 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7172 39530 7212 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7172 39450 7212 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7092 39930 7132 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7092 39850 7132 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7092 39770 7132 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7092 39690 7132 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7092 39610 7132 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7092 39530 7132 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7092 39450 7132 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7012 39930 7052 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7012 39850 7052 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7012 39770 7052 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7012 39690 7052 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7012 39610 7052 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7012 39530 7052 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 7012 39450 7052 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6932 39930 6972 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6932 39850 6972 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6932 39770 6972 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6932 39690 6972 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6932 39610 6972 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6932 39530 6972 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6932 39450 6972 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6852 39930 6892 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6852 39850 6892 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6852 39770 6892 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6852 39690 6892 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6852 39610 6892 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6852 39530 6892 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6852 39450 6892 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6772 39930 6812 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6772 39850 6812 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6772 39770 6812 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6772 39690 6812 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6772 39610 6812 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6772 39530 6812 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6772 39450 6812 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6692 39930 6732 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6692 39850 6732 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6692 39770 6732 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6692 39690 6732 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6692 39610 6732 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6692 39530 6732 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6692 39450 6732 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6612 39930 6652 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6612 39850 6652 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6612 39770 6652 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6612 39690 6652 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6612 39610 6652 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6612 39530 6652 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6612 39450 6652 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6532 39930 6572 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6532 39850 6572 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6532 39770 6572 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6532 39690 6572 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6532 39610 6572 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6532 39530 6572 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6532 39450 6572 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6452 39930 6492 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6452 39850 6492 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6452 39770 6492 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6452 39690 6492 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6452 39610 6492 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6452 39530 6492 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6452 39450 6492 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6372 39930 6412 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6372 39850 6412 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6372 39770 6412 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6372 39690 6412 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6372 39610 6412 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6372 39530 6412 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6372 39450 6412 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6292 39930 6332 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6292 39850 6332 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6292 39770 6332 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6292 39690 6332 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6292 39610 6332 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6292 39530 6332 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6292 39450 6332 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6212 39930 6252 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6212 39850 6252 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6212 39770 6252 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6212 39690 6252 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6212 39610 6252 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6212 39530 6252 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6212 39450 6252 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6132 39930 6172 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6132 39850 6172 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6132 39770 6172 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6132 39690 6172 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6132 39610 6172 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6132 39530 6172 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6132 39450 6172 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6052 39930 6092 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6052 39850 6092 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6052 39770 6092 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6052 39690 6092 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6052 39610 6092 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6052 39530 6092 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 6052 39450 6092 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5972 39930 6012 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5972 39850 6012 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5972 39770 6012 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5972 39690 6012 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5972 39610 6012 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5972 39530 6012 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5972 39450 6012 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5892 39930 5932 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5892 39850 5932 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5892 39770 5932 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5892 39690 5932 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5892 39610 5932 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5892 39530 5932 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5892 39450 5932 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5812 39930 5852 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5812 39850 5852 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5812 39770 5852 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5812 39690 5852 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5812 39610 5852 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5812 39530 5852 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5812 39450 5852 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5732 39930 5772 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5732 39850 5772 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5732 39770 5772 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5732 39690 5772 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5732 39610 5772 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5732 39530 5772 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5732 39450 5772 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5652 39930 5692 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5652 39850 5692 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5652 39770 5692 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5652 39690 5692 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5652 39610 5692 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5652 39530 5692 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5652 39450 5692 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5572 39930 5612 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5572 39850 5612 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5572 39770 5612 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5572 39690 5612 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5572 39610 5612 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5572 39530 5612 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5572 39450 5612 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5492 39930 5532 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5492 39850 5532 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5492 39770 5532 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5492 39690 5532 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5492 39610 5532 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5492 39530 5532 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5492 39450 5532 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5412 39930 5452 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5412 39850 5452 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5412 39770 5452 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5412 39690 5452 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5412 39610 5452 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5412 39530 5452 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5412 39450 5452 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5331 39930 5371 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5331 39850 5371 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5331 39770 5371 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5331 39690 5371 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5331 39610 5371 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5331 39530 5371 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5331 39450 5371 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5250 39930 5290 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5250 39850 5290 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5250 39770 5290 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5250 39690 5290 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5250 39610 5290 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5250 39530 5290 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5250 39450 5290 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5169 39930 5209 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5169 39850 5209 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5169 39770 5209 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5169 39690 5209 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5169 39610 5209 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5169 39530 5209 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5169 39450 5209 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5088 39930 5128 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5088 39850 5128 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5088 39770 5128 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5088 39690 5128 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5088 39610 5128 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5088 39530 5128 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5088 39450 5128 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5007 39930 5047 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5007 39850 5047 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5007 39770 5047 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5007 39690 5047 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5007 39610 5047 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5007 39530 5047 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 5007 39450 5047 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4926 39930 4966 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4926 39850 4966 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4926 39770 4966 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4926 39690 4966 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4926 39610 4966 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4926 39530 4966 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4926 39450 4966 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4845 39930 4885 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4845 39850 4885 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4845 39770 4885 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4845 39690 4885 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4845 39610 4885 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4845 39530 4885 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4845 39450 4885 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 6042 4861 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5956 4861 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5870 4861 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5784 4861 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5698 4861 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5612 4861 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5526 4861 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5440 4861 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5354 4861 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5268 4861 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4821 5182 4861 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4764 39930 4804 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4764 39850 4804 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4764 39770 4804 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4764 39690 4804 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4764 39610 4804 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4764 39530 4804 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4764 39450 4804 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 6042 4780 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5956 4780 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5870 4780 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5784 4780 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5698 4780 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5612 4780 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5526 4780 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5440 4780 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5354 4780 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5268 4780 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4740 5182 4780 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4683 39930 4723 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4683 39850 4723 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4683 39770 4723 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4683 39690 4723 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4683 39610 4723 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4683 39530 4723 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4683 39450 4723 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 6042 4699 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5956 4699 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5870 4699 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5784 4699 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5698 4699 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5612 4699 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5526 4699 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5440 4699 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5354 4699 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5268 4699 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4659 5182 4699 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4602 39930 4642 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4602 39850 4642 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4602 39770 4642 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4602 39690 4642 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4602 39610 4642 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4602 39530 4642 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4602 39450 4642 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 6042 4618 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5956 4618 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5870 4618 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5784 4618 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5698 4618 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5612 4618 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5526 4618 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5440 4618 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5354 4618 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5268 4618 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4578 5182 4618 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4521 39930 4561 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4521 39850 4561 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4521 39770 4561 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4521 39690 4561 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4521 39610 4561 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4521 39530 4561 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4521 39450 4561 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 6042 4537 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5956 4537 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5870 4537 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5784 4537 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5698 4537 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5612 4537 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5526 4537 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5440 4537 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5354 4537 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5268 4537 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4497 5182 4537 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4440 39930 4480 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4440 39850 4480 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4440 39770 4480 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4440 39690 4480 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4440 39610 4480 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4440 39530 4480 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4440 39450 4480 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 6042 4456 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5956 4456 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5870 4456 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5784 4456 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5698 4456 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5612 4456 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5526 4456 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5440 4456 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5354 4456 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5268 4456 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4416 5182 4456 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4359 39930 4399 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4359 39850 4399 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4359 39770 4399 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4359 39690 4399 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4359 39610 4399 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4359 39530 4399 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4359 39450 4399 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 6042 4375 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5956 4375 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5870 4375 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5784 4375 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5698 4375 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5612 4375 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5526 4375 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5440 4375 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5354 4375 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5268 4375 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4335 5182 4375 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4278 39930 4318 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4278 39850 4318 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4278 39770 4318 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4278 39690 4318 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4278 39610 4318 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4278 39530 4318 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4278 39450 4318 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 6042 4294 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5956 4294 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5870 4294 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5784 4294 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5698 4294 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5612 4294 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5526 4294 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5440 4294 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5354 4294 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5268 4294 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4254 5182 4294 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4197 39930 4237 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4197 39850 4237 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4197 39770 4237 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4197 39690 4237 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4197 39610 4237 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4197 39530 4237 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4197 39450 4237 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 6042 4213 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5956 4213 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5870 4213 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5784 4213 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5698 4213 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5612 4213 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5526 4213 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5440 4213 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5354 4213 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5268 4213 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4173 5182 4213 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4116 39930 4156 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4116 39850 4156 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4116 39770 4156 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4116 39690 4156 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4116 39610 4156 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4116 39530 4156 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4116 39450 4156 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 6042 4132 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5956 4132 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5870 4132 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5784 4132 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5698 4132 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5612 4132 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5526 4132 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5440 4132 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5354 4132 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5268 4132 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4092 5182 4132 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4035 39930 4075 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4035 39850 4075 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4035 39770 4075 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4035 39690 4075 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4035 39610 4075 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4035 39530 4075 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4035 39450 4075 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 6042 4051 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5956 4051 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5870 4051 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5784 4051 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5698 4051 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5612 4051 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5526 4051 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5440 4051 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5354 4051 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5268 4051 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 4011 5182 4051 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3954 39930 3994 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3954 39850 3994 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3954 39770 3994 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3954 39690 3994 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3954 39610 3994 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3954 39530 3994 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3954 39450 3994 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 6042 3970 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5956 3970 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5870 3970 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5784 3970 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5698 3970 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5612 3970 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5526 3970 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5440 3970 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5354 3970 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5268 3970 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3930 5182 3970 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3873 39930 3913 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3873 39850 3913 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3873 39770 3913 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3873 39690 3913 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3873 39610 3913 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3873 39530 3913 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3873 39450 3913 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 6042 3889 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5956 3889 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5870 3889 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5784 3889 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5698 3889 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5612 3889 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5526 3889 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5440 3889 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5354 3889 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5268 3889 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3849 5182 3889 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3792 39930 3832 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3792 39850 3832 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3792 39770 3832 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3792 39690 3832 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3792 39610 3832 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3792 39530 3832 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3792 39450 3832 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 6042 3808 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5956 3808 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5870 3808 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5784 3808 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5698 3808 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5612 3808 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5526 3808 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5440 3808 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5354 3808 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5268 3808 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3768 5182 3808 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3711 39930 3751 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3711 39850 3751 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3711 39770 3751 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3711 39690 3751 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3711 39610 3751 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3711 39530 3751 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3711 39450 3751 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 6042 3727 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5956 3727 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5870 3727 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5784 3727 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5698 3727 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5612 3727 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5526 3727 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5440 3727 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5354 3727 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5268 3727 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3687 5182 3727 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3630 39930 3670 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3630 39850 3670 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3630 39770 3670 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3630 39690 3670 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3630 39610 3670 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3630 39530 3670 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3630 39450 3670 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 6042 3646 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5956 3646 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5870 3646 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5784 3646 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5698 3646 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5612 3646 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5526 3646 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5440 3646 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5354 3646 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5268 3646 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3606 5182 3646 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3549 39930 3589 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3549 39850 3589 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3549 39770 3589 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3549 39690 3589 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3549 39610 3589 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3549 39530 3589 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3549 39450 3589 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 6042 3565 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5956 3565 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5870 3565 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5784 3565 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5698 3565 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5612 3565 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5526 3565 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5440 3565 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5354 3565 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5268 3565 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3525 5182 3565 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3468 39930 3508 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3468 39850 3508 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3468 39770 3508 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3468 39690 3508 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3468 39610 3508 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3468 39530 3508 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3468 39450 3508 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 6042 3484 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5956 3484 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5870 3484 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5784 3484 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5698 3484 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5612 3484 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5526 3484 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5440 3484 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5354 3484 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5268 3484 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3444 5182 3484 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3387 39930 3427 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3387 39850 3427 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3387 39770 3427 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3387 39690 3427 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3387 39610 3427 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3387 39530 3427 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3387 39450 3427 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 6042 3403 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5956 3403 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5870 3403 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5784 3403 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5698 3403 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5612 3403 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5526 3403 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5440 3403 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5354 3403 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5268 3403 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3363 5182 3403 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3306 39930 3346 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3306 39850 3346 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3306 39770 3346 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3306 39690 3346 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3306 39610 3346 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3306 39530 3346 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3306 39450 3346 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 6042 3322 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5956 3322 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5870 3322 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5784 3322 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5698 3322 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5612 3322 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5526 3322 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5440 3322 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5354 3322 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5268 3322 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3282 5182 3322 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3225 39930 3265 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3225 39850 3265 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3225 39770 3265 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3225 39690 3265 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3225 39610 3265 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3225 39530 3265 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3225 39450 3265 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 6042 3241 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5956 3241 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5870 3241 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5784 3241 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5698 3241 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5612 3241 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5526 3241 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5440 3241 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5354 3241 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5268 3241 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3201 5182 3241 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3144 39930 3184 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3144 39850 3184 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3144 39770 3184 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3144 39690 3184 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3144 39610 3184 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3144 39530 3184 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3144 39450 3184 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 6042 3160 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5956 3160 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5870 3160 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5784 3160 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5698 3160 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5612 3160 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5526 3160 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5440 3160 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5354 3160 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5268 3160 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3120 5182 3160 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3063 39930 3103 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3063 39850 3103 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3063 39770 3103 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3063 39690 3103 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3063 39610 3103 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3063 39530 3103 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3063 39450 3103 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 6042 3079 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5956 3079 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5870 3079 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5784 3079 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5698 3079 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5612 3079 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5526 3079 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5440 3079 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5354 3079 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5268 3079 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 3039 5182 3079 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2982 39930 3022 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2982 39850 3022 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2982 39770 3022 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2982 39690 3022 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2982 39610 3022 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2982 39530 3022 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2982 39450 3022 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 6042 2998 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5956 2998 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5870 2998 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5784 2998 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5698 2998 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5612 2998 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5526 2998 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5440 2998 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5354 2998 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5268 2998 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2958 5182 2998 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2901 39930 2941 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2901 39850 2941 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2901 39770 2941 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2901 39690 2941 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2901 39610 2941 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2901 39530 2941 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2901 39450 2941 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 6042 2917 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5956 2917 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5870 2917 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5784 2917 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5698 2917 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5612 2917 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5526 2917 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5440 2917 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5354 2917 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5268 2917 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2877 5182 2917 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2820 39930 2860 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2820 39850 2860 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2820 39770 2860 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2820 39690 2860 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2820 39610 2860 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2820 39530 2860 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2820 39450 2860 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 6042 2836 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5956 2836 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5870 2836 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5784 2836 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5698 2836 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5612 2836 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5526 2836 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5440 2836 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5354 2836 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5268 2836 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2796 5182 2836 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2765 39341 2805 39381 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2765 39259 2805 39299 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2739 39930 2779 39970 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2739 39850 2779 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2739 39770 2779 39810 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2739 39690 2779 39730 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2739 39610 2779 39650 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2739 39530 2779 39570 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2739 39450 2779 39490 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 6042 2755 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5956 2755 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5870 2755 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5784 2755 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5698 2755 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5612 2755 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5526 2755 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5440 2755 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5354 2755 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5268 2755 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2715 5182 2755 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 6042 2674 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5956 2674 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5870 2674 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5784 2674 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5698 2674 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5612 2674 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5526 2674 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5440 2674 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5354 2674 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5268 2674 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2634 5182 2674 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39931 2657 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39850 2657 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39769 2657 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39688 2657 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39607 2657 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39526 2657 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39445 2657 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39364 2657 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39283 2657 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39202 2657 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39121 2657 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 39040 2657 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38959 2657 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38879 2657 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38799 2657 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38719 2657 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38639 2657 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38559 2657 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38479 2657 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38399 2657 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38319 2657 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38239 2657 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38159 2657 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 38079 2657 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37999 2657 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37919 2657 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37839 2657 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37759 2657 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37679 2657 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37599 2657 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37519 2657 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37439 2657 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37359 2657 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37279 2657 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37199 2657 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37119 2657 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 37039 2657 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36959 2657 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36879 2657 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36799 2657 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36719 2657 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36639 2657 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36559 2657 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36479 2657 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36399 2657 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36319 2657 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36239 2657 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36159 2657 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 36079 2657 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35999 2657 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35919 2657 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35839 2657 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35759 2657 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35679 2657 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35599 2657 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35519 2657 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35439 2657 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35359 2657 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35279 2657 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2617 35199 2657 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 6042 2593 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5956 2593 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5870 2593 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5784 2593 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5698 2593 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5612 2593 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5526 2593 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5440 2593 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5354 2593 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5268 2593 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2553 5182 2593 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39931 2577 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39850 2577 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39769 2577 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39688 2577 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39607 2577 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39526 2577 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39445 2577 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39364 2577 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39283 2577 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39202 2577 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39121 2577 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 39040 2577 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38959 2577 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38879 2577 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38799 2577 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38719 2577 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38639 2577 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38559 2577 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38479 2577 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38399 2577 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38319 2577 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38239 2577 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38159 2577 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 38079 2577 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37999 2577 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37919 2577 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37839 2577 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37759 2577 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37679 2577 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37599 2577 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37519 2577 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37439 2577 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37359 2577 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37279 2577 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37199 2577 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37119 2577 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 37039 2577 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36959 2577 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36879 2577 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36799 2577 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36719 2577 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36639 2577 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36559 2577 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36479 2577 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36399 2577 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36319 2577 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36239 2577 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36159 2577 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 36079 2577 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35999 2577 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35919 2577 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35839 2577 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35759 2577 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35679 2577 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35599 2577 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35519 2577 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35439 2577 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35359 2577 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35279 2577 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2537 35199 2577 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 6042 2512 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5956 2512 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5870 2512 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5784 2512 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5698 2512 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5612 2512 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5526 2512 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5440 2512 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5354 2512 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5268 2512 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2472 5182 2512 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39931 2497 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39850 2497 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39769 2497 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39688 2497 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39607 2497 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39526 2497 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39445 2497 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39364 2497 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39283 2497 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39202 2497 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39121 2497 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 39040 2497 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38959 2497 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38879 2497 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38799 2497 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38719 2497 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38639 2497 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38559 2497 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38479 2497 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38399 2497 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38319 2497 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38239 2497 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38159 2497 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 38079 2497 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37999 2497 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37919 2497 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37839 2497 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37759 2497 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37679 2497 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37599 2497 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37519 2497 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37439 2497 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37359 2497 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37279 2497 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37199 2497 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37119 2497 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 37039 2497 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36959 2497 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36879 2497 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36799 2497 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36719 2497 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36639 2497 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36559 2497 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36479 2497 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36399 2497 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36319 2497 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36239 2497 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36159 2497 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 36079 2497 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35999 2497 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35919 2497 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35839 2497 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35759 2497 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35679 2497 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35599 2497 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35519 2497 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35439 2497 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35359 2497 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35279 2497 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2457 35199 2497 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 6042 2431 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5956 2431 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5870 2431 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5784 2431 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5698 2431 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5612 2431 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5526 2431 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5440 2431 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5354 2431 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5268 2431 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2391 5182 2431 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39931 2417 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39850 2417 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39769 2417 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39688 2417 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39607 2417 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39526 2417 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39445 2417 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39364 2417 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39283 2417 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39202 2417 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39121 2417 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 39040 2417 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38959 2417 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38879 2417 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38799 2417 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38719 2417 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38639 2417 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38559 2417 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38479 2417 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38399 2417 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38319 2417 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38239 2417 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38159 2417 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 38079 2417 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37999 2417 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37919 2417 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37839 2417 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37759 2417 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37679 2417 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37599 2417 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37519 2417 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37439 2417 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37359 2417 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37279 2417 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37199 2417 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37119 2417 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 37039 2417 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36959 2417 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36879 2417 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36799 2417 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36719 2417 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36639 2417 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36559 2417 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36479 2417 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36399 2417 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36319 2417 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36239 2417 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36159 2417 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 36079 2417 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35999 2417 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35919 2417 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35839 2417 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35759 2417 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35679 2417 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35599 2417 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35519 2417 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35439 2417 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35359 2417 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35279 2417 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2377 35199 2417 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 6042 2350 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5956 2350 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5870 2350 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5784 2350 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5698 2350 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5612 2350 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5526 2350 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5440 2350 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5354 2350 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5268 2350 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2310 5182 2350 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39931 2337 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39850 2337 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39769 2337 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39688 2337 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39607 2337 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39526 2337 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39445 2337 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39364 2337 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39283 2337 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39202 2337 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39121 2337 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 39040 2337 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38959 2337 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38879 2337 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38799 2337 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38719 2337 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38639 2337 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38559 2337 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38479 2337 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38399 2337 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38319 2337 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38239 2337 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38159 2337 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 38079 2337 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37999 2337 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37919 2337 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37839 2337 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37759 2337 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37679 2337 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37599 2337 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37519 2337 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37439 2337 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37359 2337 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37279 2337 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37199 2337 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37119 2337 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 37039 2337 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36959 2337 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36879 2337 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36799 2337 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36719 2337 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36639 2337 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36559 2337 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36479 2337 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36399 2337 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36319 2337 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36239 2337 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36159 2337 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 36079 2337 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35999 2337 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35919 2337 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35839 2337 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35759 2337 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35679 2337 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35599 2337 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35519 2337 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35439 2337 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35359 2337 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35279 2337 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2297 35199 2337 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 6042 2269 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5956 2269 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5870 2269 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5784 2269 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5698 2269 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5612 2269 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5526 2269 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5440 2269 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5354 2269 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5268 2269 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2229 5182 2269 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39931 2257 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39850 2257 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39769 2257 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39688 2257 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39607 2257 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39526 2257 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39445 2257 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39364 2257 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39283 2257 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39202 2257 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39121 2257 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 39040 2257 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38959 2257 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38879 2257 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38799 2257 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38719 2257 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38639 2257 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38559 2257 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38479 2257 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38399 2257 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38319 2257 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38239 2257 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38159 2257 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 38079 2257 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37999 2257 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37919 2257 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37839 2257 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37759 2257 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37679 2257 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37599 2257 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37519 2257 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37439 2257 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37359 2257 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37279 2257 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37199 2257 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37119 2257 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 37039 2257 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36959 2257 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36879 2257 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36799 2257 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36719 2257 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36639 2257 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36559 2257 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36479 2257 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36399 2257 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36319 2257 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36239 2257 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36159 2257 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 36079 2257 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35999 2257 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35919 2257 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35839 2257 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35759 2257 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35679 2257 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35599 2257 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35519 2257 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35439 2257 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35359 2257 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35279 2257 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2217 35199 2257 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 6042 2188 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5956 2188 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5870 2188 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5784 2188 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5698 2188 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5612 2188 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5526 2188 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5440 2188 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5354 2188 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5268 2188 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2148 5182 2188 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39931 2177 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39850 2177 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39769 2177 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39688 2177 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39607 2177 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39526 2177 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39445 2177 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39364 2177 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39283 2177 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39202 2177 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39121 2177 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 39040 2177 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38959 2177 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38879 2177 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38799 2177 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38719 2177 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38639 2177 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38559 2177 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38479 2177 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38399 2177 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38319 2177 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38239 2177 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38159 2177 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 38079 2177 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37999 2177 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37919 2177 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37839 2177 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37759 2177 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37679 2177 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37599 2177 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37519 2177 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37439 2177 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37359 2177 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37279 2177 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37199 2177 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37119 2177 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 37039 2177 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36959 2177 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36879 2177 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36799 2177 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36719 2177 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36639 2177 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36559 2177 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36479 2177 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36399 2177 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36319 2177 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36239 2177 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36159 2177 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 36079 2177 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35999 2177 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35919 2177 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35839 2177 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35759 2177 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35679 2177 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35599 2177 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35519 2177 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35439 2177 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35359 2177 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35279 2177 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2137 35199 2177 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 6042 2107 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5956 2107 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5870 2107 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5784 2107 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5698 2107 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5612 2107 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5526 2107 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5440 2107 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5354 2107 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5268 2107 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2067 5182 2107 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39931 2097 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39850 2097 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39769 2097 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39688 2097 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39607 2097 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39526 2097 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39445 2097 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39364 2097 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39283 2097 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39202 2097 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39121 2097 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 39040 2097 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38959 2097 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38879 2097 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38799 2097 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38719 2097 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38639 2097 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38559 2097 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38479 2097 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38399 2097 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38319 2097 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38239 2097 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38159 2097 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 38079 2097 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37999 2097 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37919 2097 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37839 2097 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37759 2097 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37679 2097 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37599 2097 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37519 2097 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37439 2097 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37359 2097 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37279 2097 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37199 2097 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37119 2097 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 37039 2097 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36959 2097 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36879 2097 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36799 2097 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36719 2097 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36639 2097 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36559 2097 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36479 2097 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36399 2097 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36319 2097 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36239 2097 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36159 2097 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 36079 2097 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35999 2097 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35919 2097 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35839 2097 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35759 2097 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35679 2097 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35599 2097 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35519 2097 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35439 2097 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35359 2097 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35279 2097 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 2057 35199 2097 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 6042 2026 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5956 2026 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5870 2026 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5784 2026 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5698 2026 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5612 2026 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5526 2026 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5440 2026 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5354 2026 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5268 2026 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1986 5182 2026 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39931 2017 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39850 2017 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39769 2017 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39688 2017 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39607 2017 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39526 2017 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39445 2017 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39364 2017 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39283 2017 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39202 2017 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39121 2017 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 39040 2017 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38959 2017 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38879 2017 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38799 2017 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38719 2017 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38639 2017 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38559 2017 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38479 2017 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38399 2017 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38319 2017 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38239 2017 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38159 2017 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 38079 2017 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37999 2017 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37919 2017 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37839 2017 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37759 2017 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37679 2017 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37599 2017 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37519 2017 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37439 2017 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37359 2017 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37279 2017 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37199 2017 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37119 2017 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 37039 2017 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36959 2017 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36879 2017 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36799 2017 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36719 2017 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36639 2017 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36559 2017 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36479 2017 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36399 2017 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36319 2017 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36239 2017 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36159 2017 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 36079 2017 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35999 2017 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35919 2017 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35839 2017 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35759 2017 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35679 2017 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35599 2017 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35519 2017 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35439 2017 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35359 2017 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35279 2017 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1977 35199 2017 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 6042 1945 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5956 1945 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5870 1945 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5784 1945 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5698 1945 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5612 1945 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5526 1945 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5440 1945 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5354 1945 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5268 1945 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1905 5182 1945 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39931 1937 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39850 1937 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39769 1937 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39688 1937 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39607 1937 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39526 1937 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39445 1937 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39364 1937 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39283 1937 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39202 1937 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39121 1937 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 39040 1937 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38959 1937 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38879 1937 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38799 1937 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38719 1937 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38639 1937 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38559 1937 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38479 1937 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38399 1937 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38319 1937 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38239 1937 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38159 1937 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 38079 1937 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37999 1937 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37919 1937 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37839 1937 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37759 1937 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37679 1937 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37599 1937 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37519 1937 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37439 1937 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37359 1937 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37279 1937 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37199 1937 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37119 1937 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 37039 1937 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36959 1937 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36879 1937 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36799 1937 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36719 1937 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36639 1937 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36559 1937 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36479 1937 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36399 1937 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36319 1937 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36239 1937 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36159 1937 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 36079 1937 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35999 1937 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35919 1937 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35839 1937 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35759 1937 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35679 1937 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35599 1937 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35519 1937 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35439 1937 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35359 1937 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35279 1937 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1897 35199 1937 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 6042 1864 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5956 1864 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5870 1864 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5784 1864 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5698 1864 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5612 1864 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5526 1864 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5440 1864 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5354 1864 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5268 1864 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1824 5182 1864 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39931 1857 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39850 1857 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39769 1857 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39688 1857 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39607 1857 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39526 1857 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39445 1857 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39364 1857 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39283 1857 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39202 1857 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39121 1857 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 39040 1857 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38959 1857 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38879 1857 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38799 1857 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38719 1857 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38639 1857 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38559 1857 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38479 1857 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38399 1857 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38319 1857 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38239 1857 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38159 1857 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 38079 1857 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37999 1857 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37919 1857 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37839 1857 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37759 1857 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37679 1857 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37599 1857 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37519 1857 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37439 1857 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37359 1857 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37279 1857 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37199 1857 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37119 1857 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 37039 1857 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36959 1857 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36879 1857 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36799 1857 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36719 1857 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36639 1857 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36559 1857 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36479 1857 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36399 1857 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36319 1857 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36239 1857 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36159 1857 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 36079 1857 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35999 1857 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35919 1857 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35839 1857 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35759 1857 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35679 1857 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35599 1857 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35519 1857 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35439 1857 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35359 1857 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35279 1857 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1817 35199 1857 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 6042 1783 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5956 1783 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5870 1783 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5784 1783 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5698 1783 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5612 1783 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5526 1783 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5440 1783 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5354 1783 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5268 1783 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1743 5182 1783 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39931 1777 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39850 1777 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39769 1777 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39688 1777 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39607 1777 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39526 1777 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39445 1777 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39364 1777 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39283 1777 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39202 1777 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39121 1777 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 39040 1777 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38959 1777 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38879 1777 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38799 1777 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38719 1777 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38639 1777 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38559 1777 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38479 1777 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38399 1777 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38319 1777 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38239 1777 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38159 1777 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 38079 1777 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37999 1777 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37919 1777 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37839 1777 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37759 1777 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37679 1777 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37599 1777 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37519 1777 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37439 1777 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37359 1777 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37279 1777 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37199 1777 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37119 1777 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 37039 1777 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36959 1777 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36879 1777 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36799 1777 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36719 1777 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36639 1777 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36559 1777 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36479 1777 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36399 1777 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36319 1777 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36239 1777 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36159 1777 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 36079 1777 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35999 1777 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35919 1777 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35839 1777 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35759 1777 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35679 1777 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35599 1777 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35519 1777 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35439 1777 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35359 1777 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35279 1777 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1737 35199 1777 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 6042 1702 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5956 1702 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5870 1702 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5784 1702 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5698 1702 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5612 1702 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5526 1702 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5440 1702 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5354 1702 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5268 1702 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1662 5182 1702 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39931 1697 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39850 1697 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39769 1697 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39688 1697 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39607 1697 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39526 1697 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39445 1697 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39364 1697 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39283 1697 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39202 1697 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39121 1697 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 39040 1697 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38959 1697 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38879 1697 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38799 1697 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38719 1697 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38639 1697 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38559 1697 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38479 1697 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38399 1697 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38319 1697 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38239 1697 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38159 1697 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 38079 1697 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37999 1697 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37919 1697 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37839 1697 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37759 1697 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37679 1697 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37599 1697 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37519 1697 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37439 1697 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37359 1697 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37279 1697 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37199 1697 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37119 1697 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 37039 1697 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36959 1697 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36879 1697 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36799 1697 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36719 1697 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36639 1697 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36559 1697 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36479 1697 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36399 1697 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36319 1697 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36239 1697 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36159 1697 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 36079 1697 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35999 1697 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35919 1697 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35839 1697 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35759 1697 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35679 1697 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35599 1697 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35519 1697 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35439 1697 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35359 1697 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35279 1697 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1657 35199 1697 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 6042 1621 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5956 1621 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5870 1621 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5784 1621 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5698 1621 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5612 1621 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5526 1621 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5440 1621 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5354 1621 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5268 1621 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1581 5182 1621 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39931 1617 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39850 1617 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39769 1617 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39688 1617 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39607 1617 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39526 1617 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39445 1617 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39364 1617 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39283 1617 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39202 1617 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39121 1617 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 39040 1617 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38959 1617 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38879 1617 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38799 1617 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38719 1617 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38639 1617 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38559 1617 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38479 1617 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38399 1617 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38319 1617 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38239 1617 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38159 1617 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 38079 1617 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37999 1617 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37919 1617 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37839 1617 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37759 1617 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37679 1617 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37599 1617 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37519 1617 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37439 1617 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37359 1617 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37279 1617 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37199 1617 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37119 1617 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 37039 1617 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36959 1617 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36879 1617 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36799 1617 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36719 1617 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36639 1617 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36559 1617 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36479 1617 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36399 1617 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36319 1617 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36239 1617 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36159 1617 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 36079 1617 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35999 1617 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35919 1617 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35839 1617 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35759 1617 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35679 1617 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35599 1617 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35519 1617 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35439 1617 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35359 1617 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35279 1617 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1577 35199 1617 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 6042 1540 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5956 1540 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5870 1540 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5784 1540 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5698 1540 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5612 1540 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5526 1540 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5440 1540 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5354 1540 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5268 1540 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1500 5182 1540 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39931 1537 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39850 1537 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39769 1537 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39688 1537 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39607 1537 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39526 1537 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39445 1537 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39364 1537 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39283 1537 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39202 1537 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39121 1537 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 39040 1537 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38959 1537 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38879 1537 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38799 1537 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38719 1537 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38639 1537 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38559 1537 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38479 1537 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38399 1537 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38319 1537 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38239 1537 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38159 1537 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 38079 1537 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37999 1537 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37919 1537 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37839 1537 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37759 1537 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37679 1537 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37599 1537 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37519 1537 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37439 1537 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37359 1537 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37279 1537 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37199 1537 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37119 1537 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 37039 1537 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36959 1537 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36879 1537 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36799 1537 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36719 1537 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36639 1537 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36559 1537 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36479 1537 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36399 1537 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36319 1537 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36239 1537 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36159 1537 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 36079 1537 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35999 1537 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35919 1537 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35839 1537 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35759 1537 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35679 1537 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35599 1537 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35519 1537 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35439 1537 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35359 1537 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35279 1537 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1497 35199 1537 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 6042 1459 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5956 1459 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5870 1459 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5784 1459 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5698 1459 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5612 1459 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5526 1459 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5440 1459 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5354 1459 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5268 1459 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1419 5182 1459 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39931 1457 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39850 1457 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39769 1457 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39688 1457 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39607 1457 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39526 1457 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39445 1457 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39364 1457 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39283 1457 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39202 1457 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39121 1457 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 39040 1457 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38959 1457 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38879 1457 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38799 1457 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38719 1457 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38639 1457 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38559 1457 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38479 1457 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38399 1457 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38319 1457 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38239 1457 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38159 1457 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 38079 1457 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37999 1457 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37919 1457 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37839 1457 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37759 1457 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37679 1457 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37599 1457 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37519 1457 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37439 1457 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37359 1457 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37279 1457 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37199 1457 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37119 1457 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 37039 1457 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36959 1457 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36879 1457 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36799 1457 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36719 1457 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36639 1457 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36559 1457 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36479 1457 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36399 1457 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36319 1457 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36239 1457 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36159 1457 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 36079 1457 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35999 1457 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35919 1457 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35839 1457 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35759 1457 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35679 1457 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35599 1457 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35519 1457 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35439 1457 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35359 1457 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35279 1457 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1417 35199 1457 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 6042 1378 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5956 1378 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5870 1378 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5784 1378 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5698 1378 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5612 1378 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5526 1378 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5440 1378 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5354 1378 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5268 1378 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1338 5182 1378 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39931 1377 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39850 1377 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39769 1377 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39688 1377 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39607 1377 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39526 1377 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39445 1377 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39364 1377 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39283 1377 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39202 1377 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39121 1377 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 39040 1377 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38959 1377 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38879 1377 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38799 1377 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38719 1377 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38639 1377 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38559 1377 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38479 1377 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38399 1377 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38319 1377 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38239 1377 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38159 1377 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 38079 1377 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37999 1377 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37919 1377 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37839 1377 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37759 1377 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37679 1377 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37599 1377 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37519 1377 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37439 1377 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37359 1377 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37279 1377 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37199 1377 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37119 1377 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 37039 1377 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36959 1377 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36879 1377 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36799 1377 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36719 1377 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36639 1377 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36559 1377 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36479 1377 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36399 1377 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36319 1377 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36239 1377 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36159 1377 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 36079 1377 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35999 1377 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35919 1377 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35839 1377 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35759 1377 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35679 1377 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35599 1377 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35519 1377 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35439 1377 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35359 1377 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35279 1377 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1337 35199 1377 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39931 1297 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39850 1297 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39769 1297 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39688 1297 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39607 1297 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39526 1297 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39445 1297 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39364 1297 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39283 1297 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39202 1297 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39121 1297 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 39040 1297 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38959 1297 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38879 1297 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38799 1297 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38719 1297 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38639 1297 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38559 1297 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38479 1297 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38399 1297 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38319 1297 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38239 1297 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38159 1297 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 38079 1297 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37999 1297 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37919 1297 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37839 1297 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37759 1297 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37679 1297 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37599 1297 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37519 1297 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37439 1297 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37359 1297 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37279 1297 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37199 1297 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37119 1297 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 37039 1297 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36959 1297 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36879 1297 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36799 1297 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36719 1297 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36639 1297 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36559 1297 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36479 1297 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36399 1297 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36319 1297 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36239 1297 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36159 1297 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 36079 1297 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35999 1297 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35919 1297 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35839 1297 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35759 1297 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35679 1297 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35599 1297 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35519 1297 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35439 1297 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35359 1297 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35279 1297 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 35199 1297 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 6042 1297 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5956 1297 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5870 1297 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5784 1297 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5698 1297 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5612 1297 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5526 1297 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5440 1297 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5354 1297 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5268 1297 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1257 5182 1297 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39931 1217 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39850 1217 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39769 1217 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39688 1217 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39607 1217 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39526 1217 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39445 1217 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39364 1217 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39283 1217 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39202 1217 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39121 1217 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 39040 1217 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38959 1217 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38879 1217 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38799 1217 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38719 1217 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38639 1217 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38559 1217 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38479 1217 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38399 1217 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38319 1217 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38239 1217 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38159 1217 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 38079 1217 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37999 1217 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37919 1217 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37839 1217 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37759 1217 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37679 1217 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37599 1217 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37519 1217 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37439 1217 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37359 1217 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37279 1217 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37199 1217 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37119 1217 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 37039 1217 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36959 1217 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36879 1217 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36799 1217 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36719 1217 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36639 1217 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36559 1217 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36479 1217 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36399 1217 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36319 1217 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36239 1217 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36159 1217 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 36079 1217 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35999 1217 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35919 1217 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35839 1217 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35759 1217 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35679 1217 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35599 1217 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35519 1217 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35439 1217 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35359 1217 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35279 1217 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1177 35199 1217 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 6042 1216 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5956 1216 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5870 1216 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5784 1216 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5698 1216 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5612 1216 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5526 1216 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5440 1216 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5354 1216 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5268 1216 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1176 5182 1216 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39931 1137 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39850 1137 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39769 1137 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39688 1137 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39607 1137 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39526 1137 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39445 1137 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39364 1137 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39283 1137 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39202 1137 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39121 1137 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 39040 1137 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38959 1137 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38879 1137 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38799 1137 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38719 1137 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38639 1137 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38559 1137 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38479 1137 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38399 1137 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38319 1137 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38239 1137 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38159 1137 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 38079 1137 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37999 1137 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37919 1137 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37839 1137 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37759 1137 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37679 1137 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37599 1137 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37519 1137 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37439 1137 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37359 1137 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37279 1137 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37199 1137 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37119 1137 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 37039 1137 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36959 1137 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36879 1137 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36799 1137 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36719 1137 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36639 1137 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36559 1137 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36479 1137 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36399 1137 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36319 1137 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36239 1137 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36159 1137 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 36079 1137 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35999 1137 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35919 1137 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35839 1137 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35759 1137 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35679 1137 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35599 1137 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35519 1137 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35439 1137 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35359 1137 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35279 1137 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1097 35199 1137 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 6042 1135 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5956 1135 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5870 1135 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5784 1135 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5698 1135 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5612 1135 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5526 1135 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5440 1135 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5354 1135 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5268 1135 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1095 5182 1135 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39931 1057 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39850 1057 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39769 1057 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39688 1057 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39607 1057 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39526 1057 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39445 1057 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39364 1057 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39283 1057 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39202 1057 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39121 1057 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 39040 1057 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38959 1057 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38879 1057 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38799 1057 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38719 1057 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38639 1057 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38559 1057 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38479 1057 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38399 1057 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38319 1057 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38239 1057 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38159 1057 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 38079 1057 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37999 1057 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37919 1057 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37839 1057 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37759 1057 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37679 1057 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37599 1057 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37519 1057 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37439 1057 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37359 1057 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37279 1057 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37199 1057 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37119 1057 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 37039 1057 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36959 1057 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36879 1057 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36799 1057 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36719 1057 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36639 1057 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36559 1057 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36479 1057 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36399 1057 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36319 1057 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36239 1057 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36159 1057 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 36079 1057 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35999 1057 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35919 1057 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35839 1057 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35759 1057 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35679 1057 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35599 1057 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35519 1057 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35439 1057 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35359 1057 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35279 1057 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1017 35199 1057 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 6042 1054 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5956 1054 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5870 1054 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5784 1054 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5698 1054 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5612 1054 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5526 1054 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5440 1054 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5354 1054 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5268 1054 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 1014 5182 1054 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39931 977 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39850 977 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39769 977 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39688 977 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39607 977 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39526 977 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39445 977 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39364 977 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39283 977 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39202 977 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39121 977 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 39040 977 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38959 977 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38879 977 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38799 977 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38719 977 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38639 977 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38559 977 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38479 977 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38399 977 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38319 977 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38239 977 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38159 977 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 38079 977 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37999 977 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37919 977 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37839 977 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37759 977 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37679 977 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37599 977 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37519 977 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37439 977 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37359 977 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37279 977 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37199 977 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37119 977 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 37039 977 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36959 977 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36879 977 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36799 977 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36719 977 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36639 977 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36559 977 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36479 977 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36399 977 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36319 977 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36239 977 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36159 977 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 36079 977 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35999 977 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35919 977 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35839 977 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35759 977 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35679 977 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35599 977 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35519 977 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35439 977 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35359 977 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35279 977 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 937 35199 977 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 6042 973 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5956 973 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5870 973 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5784 973 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5698 973 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5612 973 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5526 973 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5440 973 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5354 973 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5268 973 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 933 5182 973 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39931 897 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39850 897 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39769 897 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39688 897 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39607 897 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39526 897 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39445 897 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39364 897 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39283 897 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39202 897 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39121 897 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 39040 897 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38959 897 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38879 897 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38799 897 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38719 897 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38639 897 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38559 897 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38479 897 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38399 897 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38319 897 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38239 897 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38159 897 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 38079 897 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37999 897 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37919 897 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37839 897 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37759 897 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37679 897 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37599 897 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37519 897 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37439 897 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37359 897 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37279 897 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37199 897 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37119 897 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 37039 897 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36959 897 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36879 897 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36799 897 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36719 897 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36639 897 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36559 897 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36479 897 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36399 897 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36319 897 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36239 897 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36159 897 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 36079 897 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35999 897 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35919 897 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35839 897 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35759 897 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35679 897 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35599 897 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35519 897 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35439 897 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35359 897 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35279 897 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 857 35199 897 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 6042 892 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5956 892 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5870 892 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5784 892 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5698 892 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5612 892 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5526 892 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5440 892 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5354 892 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5268 892 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 852 5182 892 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39931 817 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39850 817 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39769 817 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39688 817 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39607 817 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39526 817 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39445 817 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39364 817 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39283 817 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39202 817 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39121 817 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 39040 817 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38959 817 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38879 817 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38799 817 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38719 817 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38639 817 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38559 817 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38479 817 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38399 817 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38319 817 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38239 817 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38159 817 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 38079 817 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37999 817 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37919 817 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37839 817 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37759 817 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37679 817 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37599 817 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37519 817 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37439 817 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37359 817 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37279 817 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37199 817 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37119 817 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 37039 817 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36959 817 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36879 817 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36799 817 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36719 817 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36639 817 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36559 817 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36479 817 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36399 817 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36319 817 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36239 817 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36159 817 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 36079 817 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35999 817 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35919 817 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35839 817 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35759 817 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35679 817 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35599 817 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35519 817 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35439 817 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35359 817 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35279 817 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 777 35199 817 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 6042 811 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5956 811 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5870 811 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5784 811 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5698 811 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5612 811 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5526 811 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5440 811 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5354 811 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5268 811 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 771 5182 811 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39931 737 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39850 737 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39769 737 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39688 737 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39607 737 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39526 737 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39445 737 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39364 737 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39283 737 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39202 737 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39121 737 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 39040 737 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38959 737 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38879 737 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38799 737 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38719 737 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38639 737 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38559 737 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38479 737 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38399 737 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38319 737 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38239 737 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38159 737 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 38079 737 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37999 737 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37919 737 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37839 737 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37759 737 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37679 737 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37599 737 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37519 737 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37439 737 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37359 737 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37279 737 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37199 737 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37119 737 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 37039 737 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36959 737 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36879 737 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36799 737 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36719 737 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36639 737 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36559 737 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36479 737 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36399 737 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36319 737 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36239 737 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36159 737 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 36079 737 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35999 737 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35919 737 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35839 737 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35759 737 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35679 737 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35599 737 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35519 737 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35439 737 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35359 737 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35279 737 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 697 35199 737 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 6042 730 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5956 730 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5870 730 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5784 730 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5698 730 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5612 730 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5526 730 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5440 730 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5354 730 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5268 730 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 690 5182 730 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39931 657 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39850 657 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39769 657 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39688 657 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39607 657 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39526 657 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39445 657 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39364 657 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39283 657 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39202 657 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39121 657 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 39040 657 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38959 657 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38879 657 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38799 657 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38719 657 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38639 657 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38559 657 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38479 657 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38399 657 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38319 657 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38239 657 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38159 657 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 38079 657 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37999 657 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37919 657 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37839 657 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37759 657 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37679 657 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37599 657 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37519 657 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37439 657 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37359 657 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37279 657 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37199 657 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37119 657 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 37039 657 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36959 657 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36879 657 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36799 657 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36719 657 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36639 657 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36559 657 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36479 657 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36399 657 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36319 657 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36239 657 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36159 657 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 36079 657 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35999 657 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35919 657 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35839 657 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35759 657 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35679 657 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35599 657 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35519 657 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35439 657 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35359 657 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35279 657 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 617 35199 657 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 6042 649 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5956 649 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5870 649 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5784 649 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5698 649 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5612 649 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5526 649 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5440 649 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5354 649 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5268 649 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 609 5182 649 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39931 577 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39850 577 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39769 577 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39688 577 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39607 577 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39526 577 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39445 577 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39364 577 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39283 577 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39202 577 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39121 577 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 39040 577 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38959 577 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38879 577 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38799 577 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38719 577 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38639 577 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38559 577 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38479 577 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38399 577 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38319 577 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38239 577 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38159 577 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 38079 577 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37999 577 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37919 577 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37839 577 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37759 577 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37679 577 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37599 577 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37519 577 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37439 577 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37359 577 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37279 577 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37199 577 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37119 577 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 37039 577 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36959 577 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36879 577 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36799 577 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36719 577 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36639 577 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36559 577 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36479 577 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36399 577 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36319 577 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36239 577 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36159 577 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 36079 577 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35999 577 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35919 577 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35839 577 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35759 577 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35679 577 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35599 577 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35519 577 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35439 577 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35359 577 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35279 577 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 537 35199 577 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 6042 567 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5956 567 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5870 567 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5784 567 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5698 567 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5612 567 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5526 567 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5440 567 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5354 567 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5268 567 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 527 5182 567 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39931 497 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39850 497 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39769 497 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39688 497 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39607 497 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39526 497 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39445 497 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39364 497 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39283 497 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39202 497 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39121 497 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 39040 497 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38959 497 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38879 497 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38799 497 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38719 497 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38639 497 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38559 497 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38479 497 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38399 497 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38319 497 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38239 497 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38159 497 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 38079 497 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37999 497 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37919 497 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37839 497 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37759 497 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37679 497 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37599 497 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37519 497 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37439 497 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37359 497 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37279 497 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37199 497 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37119 497 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 37039 497 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36959 497 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36879 497 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36799 497 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36719 497 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36639 497 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36559 497 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36479 497 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36399 497 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36319 497 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36239 497 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36159 497 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 36079 497 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35999 497 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35919 497 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35839 497 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35759 497 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35679 497 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35599 497 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35519 497 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35439 497 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35359 497 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35279 497 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 457 35199 497 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 6042 485 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5956 485 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5870 485 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5784 485 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5698 485 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5612 485 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5526 485 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5440 485 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5354 485 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5268 485 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 445 5182 485 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39931 417 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39850 417 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39769 417 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39688 417 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39607 417 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39526 417 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39445 417 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39364 417 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39283 417 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39202 417 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39121 417 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 39040 417 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38959 417 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38879 417 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38799 417 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38719 417 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38639 417 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38559 417 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38479 417 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38399 417 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38319 417 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38239 417 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38159 417 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 38079 417 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37999 417 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37919 417 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37839 417 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37759 417 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37679 417 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37599 417 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37519 417 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37439 417 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37359 417 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37279 417 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37199 417 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37119 417 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 37039 417 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36959 417 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36879 417 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36799 417 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36719 417 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36639 417 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36559 417 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36479 417 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36399 417 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36319 417 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36239 417 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36159 417 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 36079 417 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35999 417 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35919 417 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35839 417 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35759 417 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35679 417 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35599 417 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35519 417 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35439 417 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35359 417 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35279 417 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 377 35199 417 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 6042 403 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5956 403 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5870 403 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5784 403 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5698 403 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5612 403 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5526 403 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5440 403 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5354 403 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5268 403 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 363 5182 403 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39931 337 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39850 337 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39769 337 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39688 337 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39607 337 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39526 337 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39445 337 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39364 337 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39283 337 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39202 337 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39121 337 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 39040 337 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38959 337 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38879 337 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38799 337 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38719 337 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38639 337 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38559 337 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38479 337 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38399 337 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38319 337 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38239 337 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38159 337 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 38079 337 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37999 337 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37919 337 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37839 337 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37759 337 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37679 337 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37599 337 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37519 337 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37439 337 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37359 337 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37279 337 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37199 337 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37119 337 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 37039 337 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36959 337 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36879 337 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36799 337 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36719 337 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36639 337 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36559 337 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36479 337 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36399 337 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36319 337 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36239 337 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36159 337 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 36079 337 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35999 337 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35919 337 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35839 337 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35759 337 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35679 337 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35599 337 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35519 337 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35439 337 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35359 337 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35279 337 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 297 35199 337 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 6042 321 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5956 321 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5870 321 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5784 321 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5698 321 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5612 321 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5526 321 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5440 321 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5354 321 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5268 321 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 281 5182 321 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39931 257 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39850 257 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39769 257 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39688 257 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39607 257 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39526 257 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39445 257 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39364 257 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39283 257 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39202 257 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39121 257 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 39040 257 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38959 257 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38879 257 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38799 257 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38719 257 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38639 257 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38559 257 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38479 257 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38399 257 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38319 257 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38239 257 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38159 257 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 38079 257 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37999 257 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37919 257 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37839 257 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37759 257 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37679 257 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37599 257 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37519 257 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37439 257 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37359 257 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37279 257 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37199 257 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37119 257 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 37039 257 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36959 257 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36879 257 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36799 257 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36719 257 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36639 257 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36559 257 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36479 257 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36399 257 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36319 257 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36239 257 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36159 257 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 36079 257 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35999 257 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35919 257 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35839 257 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35759 257 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35679 257 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35599 257 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35519 257 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35439 257 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35359 257 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35279 257 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 217 35199 257 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 6042 239 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5956 239 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5870 239 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5784 239 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5698 239 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5612 239 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5526 239 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5440 239 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5354 239 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5268 239 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 199 5182 239 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39931 177 39971 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39850 177 39890 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39769 177 39809 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39688 177 39728 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39607 177 39647 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39526 177 39566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39445 177 39485 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39364 177 39404 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39283 177 39323 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39202 177 39242 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39121 177 39161 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 39040 177 39080 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38959 177 38999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38879 177 38919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38799 177 38839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38719 177 38759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38639 177 38679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38559 177 38599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38479 177 38519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38399 177 38439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38319 177 38359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38239 177 38279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38159 177 38199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 38079 177 38119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37999 177 38039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37919 177 37959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37839 177 37879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37759 177 37799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37679 177 37719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37599 177 37639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37519 177 37559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37439 177 37479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37359 177 37399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37279 177 37319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37199 177 37239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37119 177 37159 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 37039 177 37079 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36959 177 36999 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36879 177 36919 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36799 177 36839 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36719 177 36759 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36639 177 36679 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36559 177 36599 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36479 177 36519 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36399 177 36439 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36319 177 36359 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36239 177 36279 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36159 177 36199 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 36079 177 36119 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35999 177 36039 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35919 177 35959 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35839 177 35879 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35759 177 35799 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35679 177 35719 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35599 177 35639 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35519 177 35559 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35439 177 35479 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35359 177 35399 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35279 177 35319 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 137 35199 177 35239 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 6042 157 6082 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5956 157 5996 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5870 157 5910 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5784 157 5824 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5698 157 5738 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5612 157 5652 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5526 157 5566 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5440 157 5480 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5354 157 5394 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5268 157 5308 1 VSSIO
port 51 nsew ground bidirectional
rlabel via3 s 117 5182 157 5222 1 VSSIO
port 51 nsew ground bidirectional
rlabel metal3 s 10078 11648 14858 12536 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal4 s 0 11647 4874 12537 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal4 s 10083 11647 15000 12537 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 12482 14840 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 12400 14840 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 12318 14840 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 12236 14840 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 12154 14840 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 12072 14840 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 11990 14840 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 11908 14840 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 11826 14840 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 11744 14840 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14800 11662 14840 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 12482 14759 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 12400 14759 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 12318 14759 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 12236 14759 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 12154 14759 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 12072 14759 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 11990 14759 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 11908 14759 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 11826 14759 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 11744 14759 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14719 11662 14759 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 12482 14678 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 12400 14678 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 12318 14678 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 12236 14678 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 12154 14678 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 12072 14678 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 11990 14678 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 11908 14678 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 11826 14678 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 11744 14678 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14638 11662 14678 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 12482 14597 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 12400 14597 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 12318 14597 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 12236 14597 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 12154 14597 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 12072 14597 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 11990 14597 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 11908 14597 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 11826 14597 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 11744 14597 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14557 11662 14597 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 12482 14516 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 12400 14516 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 12318 14516 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 12236 14516 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 12154 14516 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 12072 14516 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 11990 14516 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 11908 14516 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 11826 14516 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 11744 14516 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14476 11662 14516 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 12482 14435 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 12400 14435 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 12318 14435 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 12236 14435 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 12154 14435 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 12072 14435 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 11990 14435 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 11908 14435 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 11826 14435 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 11744 14435 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14395 11662 14435 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 12482 14354 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 12400 14354 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 12318 14354 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 12236 14354 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 12154 14354 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 12072 14354 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 11990 14354 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 11908 14354 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 11826 14354 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 11744 14354 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14314 11662 14354 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 12482 14273 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 12400 14273 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 12318 14273 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 12236 14273 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 12154 14273 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 12072 14273 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 11990 14273 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 11908 14273 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 11826 14273 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 11744 14273 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14233 11662 14273 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 12482 14192 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 12400 14192 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 12318 14192 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 12236 14192 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 12154 14192 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 12072 14192 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 11990 14192 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 11908 14192 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 11826 14192 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 11744 14192 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14152 11662 14192 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 12482 14111 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 12400 14111 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 12318 14111 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 12236 14111 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 12154 14111 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 12072 14111 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 11990 14111 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 11908 14111 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 11826 14111 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 11744 14111 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 14071 11662 14111 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 12482 14030 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 12400 14030 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 12318 14030 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 12236 14030 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 12154 14030 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 12072 14030 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 11990 14030 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 11908 14030 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 11826 14030 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 11744 14030 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13990 11662 14030 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 12482 13949 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 12400 13949 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 12318 13949 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 12236 13949 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 12154 13949 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 12072 13949 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 11990 13949 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 11908 13949 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 11826 13949 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 11744 13949 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13909 11662 13949 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 12482 13868 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 12400 13868 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 12318 13868 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 12236 13868 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 12154 13868 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 12072 13868 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 11990 13868 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 11908 13868 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 11826 13868 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 11744 13868 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13828 11662 13868 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 12482 13787 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 12400 13787 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 12318 13787 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 12236 13787 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 12154 13787 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 12072 13787 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 11990 13787 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 11908 13787 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 11826 13787 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 11744 13787 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13747 11662 13787 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 12482 13706 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 12400 13706 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 12318 13706 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 12236 13706 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 12154 13706 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 12072 13706 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 11990 13706 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 11908 13706 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 11826 13706 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 11744 13706 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13666 11662 13706 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 12482 13625 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 12400 13625 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 12318 13625 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 12236 13625 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 12154 13625 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 12072 13625 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 11990 13625 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 11908 13625 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 11826 13625 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 11744 13625 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13585 11662 13625 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 12482 13544 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 12400 13544 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 12318 13544 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 12236 13544 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 12154 13544 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 12072 13544 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 11990 13544 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 11908 13544 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 11826 13544 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 11744 13544 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13504 11662 13544 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 12482 13463 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 12400 13463 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 12318 13463 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 12236 13463 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 12154 13463 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 12072 13463 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 11990 13463 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 11908 13463 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 11826 13463 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 11744 13463 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13423 11662 13463 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 12482 13382 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 12400 13382 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 12318 13382 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 12236 13382 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 12154 13382 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 12072 13382 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 11990 13382 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 11908 13382 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 11826 13382 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 11744 13382 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13342 11662 13382 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 12482 13301 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 12400 13301 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 12318 13301 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 12236 13301 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 12154 13301 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 12072 13301 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 11990 13301 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 11908 13301 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 11826 13301 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 11744 13301 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13261 11662 13301 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 12482 13220 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 12400 13220 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 12318 13220 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 12236 13220 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 12154 13220 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 12072 13220 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 11990 13220 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 11908 13220 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 11826 13220 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 11744 13220 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13180 11662 13220 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 12482 13139 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 12400 13139 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 12318 13139 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 12236 13139 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 12154 13139 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 12072 13139 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 11990 13139 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 11908 13139 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 11826 13139 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 11744 13139 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13099 11662 13139 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 12482 13058 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 12400 13058 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 12318 13058 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 12236 13058 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 12154 13058 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 12072 13058 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 11990 13058 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 11908 13058 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 11826 13058 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 11744 13058 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 13018 11662 13058 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 12482 12977 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 12400 12977 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 12318 12977 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 12236 12977 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 12154 12977 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 12072 12977 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 11990 12977 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 11908 12977 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 11826 12977 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 11744 12977 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12937 11662 12977 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 12482 12896 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 12400 12896 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 12318 12896 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 12236 12896 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 12154 12896 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 12072 12896 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 11990 12896 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 11908 12896 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 11826 12896 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 11744 12896 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12856 11662 12896 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 12482 12815 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 12400 12815 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 12318 12815 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 12236 12815 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 12154 12815 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 12072 12815 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 11990 12815 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 11908 12815 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 11826 12815 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 11744 12815 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12775 11662 12815 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 12482 12734 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 12400 12734 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 12318 12734 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 12236 12734 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 12154 12734 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 12072 12734 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 11990 12734 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 11908 12734 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 11826 12734 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 11744 12734 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12694 11662 12734 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 12482 12653 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 12400 12653 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 12318 12653 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 12236 12653 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 12154 12653 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 12072 12653 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 11990 12653 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 11908 12653 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 11826 12653 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 11744 12653 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12613 11662 12653 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 12482 12572 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 12400 12572 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 12318 12572 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 12236 12572 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 12154 12572 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 12072 12572 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 11990 12572 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 11908 12572 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 11826 12572 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 11744 12572 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12532 11662 12572 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 12482 12491 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 12400 12491 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 12318 12491 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 12236 12491 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 12154 12491 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 12072 12491 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 11990 12491 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 11908 12491 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 11826 12491 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 11744 12491 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12451 11662 12491 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 12482 12410 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 12400 12410 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 12318 12410 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 12236 12410 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 12154 12410 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 12072 12410 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 11990 12410 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 11908 12410 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 11826 12410 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 11744 12410 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12370 11662 12410 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 12482 12329 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 12400 12329 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 12318 12329 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 12236 12329 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 12154 12329 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 12072 12329 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 11990 12329 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 11908 12329 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 11826 12329 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 11744 12329 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12289 11662 12329 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 12482 12248 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 12400 12248 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 12318 12248 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 12236 12248 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 12154 12248 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 12072 12248 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 11990 12248 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 11908 12248 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 11826 12248 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 11744 12248 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12208 11662 12248 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 12482 12167 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 12400 12167 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 12318 12167 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 12236 12167 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 12154 12167 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 12072 12167 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 11990 12167 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 11908 12167 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 11826 12167 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 11744 12167 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12127 11662 12167 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 12482 12086 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 12400 12086 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 12318 12086 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 12236 12086 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 12154 12086 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 12072 12086 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 11990 12086 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 11908 12086 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 11826 12086 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 11744 12086 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 12046 11662 12086 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 12482 12005 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 12400 12005 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 12318 12005 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 12236 12005 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 12154 12005 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 12072 12005 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 11990 12005 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 11908 12005 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 11826 12005 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 11744 12005 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11965 11662 12005 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 12482 11924 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 12400 11924 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 12318 11924 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 12236 11924 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 12154 11924 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 12072 11924 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 11990 11924 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 11908 11924 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 11826 11924 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 11744 11924 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11884 11662 11924 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 12482 11843 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 12400 11843 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 12318 11843 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 12236 11843 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 12154 11843 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 12072 11843 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 11990 11843 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 11908 11843 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 11826 11843 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 11744 11843 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11803 11662 11843 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 12482 11762 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 12400 11762 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 12318 11762 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 12236 11762 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 12154 11762 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 12072 11762 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 11990 11762 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 11908 11762 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 11826 11762 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 11744 11762 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11722 11662 11762 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 12482 11681 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 12400 11681 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 12318 11681 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 12236 11681 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 12154 11681 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 12072 11681 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 11990 11681 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 11908 11681 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 11826 11681 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 11744 11681 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11641 11662 11681 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 12482 11600 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 12400 11600 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 12318 11600 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 12236 11600 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 12154 11600 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 12072 11600 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 11990 11600 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 11908 11600 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 11826 11600 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 11744 11600 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11560 11662 11600 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 12482 11519 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 12400 11519 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 12318 11519 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 12236 11519 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 12154 11519 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 12072 11519 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 11990 11519 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 11908 11519 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 11826 11519 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 11744 11519 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11479 11662 11519 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 12482 11438 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 12400 11438 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 12318 11438 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 12236 11438 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 12154 11438 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 12072 11438 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 11990 11438 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 11908 11438 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 11826 11438 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 11744 11438 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11398 11662 11438 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 12482 11357 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 12400 11357 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 12318 11357 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 12236 11357 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 12154 11357 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 12072 11357 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 11990 11357 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 11908 11357 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 11826 11357 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 11744 11357 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11317 11662 11357 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 12482 11276 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 12400 11276 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 12318 11276 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 12236 11276 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 12154 11276 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 12072 11276 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 11990 11276 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 11908 11276 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 11826 11276 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 11744 11276 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11236 11662 11276 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 12482 11195 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 12400 11195 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 12318 11195 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 12236 11195 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 12154 11195 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 12072 11195 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 11990 11195 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 11908 11195 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 11826 11195 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 11744 11195 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11155 11662 11195 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 12482 11114 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 12400 11114 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 12318 11114 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 12236 11114 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 12154 11114 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 12072 11114 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 11990 11114 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 11908 11114 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 11826 11114 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 11744 11114 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 11074 11662 11114 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 12482 11033 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 12400 11033 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 12318 11033 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 12236 11033 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 12154 11033 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 12072 11033 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 11990 11033 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 11908 11033 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 11826 11033 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 11744 11033 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10993 11662 11033 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 12482 10952 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 12400 10952 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 12318 10952 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 12236 10952 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 12154 10952 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 12072 10952 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 11990 10952 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 11908 10952 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 11826 10952 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 11744 10952 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10912 11662 10952 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 12482 10871 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 12400 10871 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 12318 10871 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 12236 10871 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 12154 10871 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 12072 10871 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 11990 10871 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 11908 10871 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 11826 10871 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 11744 10871 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10831 11662 10871 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 12482 10790 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 12400 10790 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 12318 10790 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 12236 10790 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 12154 10790 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 12072 10790 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 11990 10790 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 11908 10790 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 11826 10790 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 11744 10790 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10750 11662 10790 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 12482 10709 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 12400 10709 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 12318 10709 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 12236 10709 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 12154 10709 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 12072 10709 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 11990 10709 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 11908 10709 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 11826 10709 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 11744 10709 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10669 11662 10709 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 12482 10628 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 12400 10628 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 12318 10628 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 12236 10628 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 12154 10628 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 12072 10628 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 11990 10628 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 11908 10628 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 11826 10628 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 11744 10628 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10588 11662 10628 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 12482 10546 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 12400 10546 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 12318 10546 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 12236 10546 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 12154 10546 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 12072 10546 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 11990 10546 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 11908 10546 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 11826 10546 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 11744 10546 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10506 11662 10546 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 12482 10464 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 12400 10464 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 12318 10464 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 12236 10464 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 12154 10464 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 12072 10464 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 11990 10464 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 11908 10464 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 11826 10464 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 11744 10464 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10424 11662 10464 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 12482 10382 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 12400 10382 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 12318 10382 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 12236 10382 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 12154 10382 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 12072 10382 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 11990 10382 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 11908 10382 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 11826 10382 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 11744 10382 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10342 11662 10382 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 12482 10300 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 12400 10300 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 12318 10300 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 12236 10300 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 12154 10300 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 12072 10300 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 11990 10300 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 11908 10300 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 11826 10300 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 11744 10300 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10260 11662 10300 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 12482 10218 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 12400 10218 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 12318 10218 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 12236 10218 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 12154 10218 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 12072 10218 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 11990 10218 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 11908 10218 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 11826 10218 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 11744 10218 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10178 11662 10218 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 12482 10136 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 12400 10136 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 12318 10136 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 12236 10136 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 12154 10136 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 12072 10136 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 11990 10136 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 11908 10136 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 11826 10136 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 11744 10136 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 10096 11662 10136 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 12482 4861 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 12400 4861 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 12318 4861 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 12236 4861 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 12154 4861 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 12072 4861 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 11990 4861 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 11908 4861 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 11826 4861 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 11744 4861 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4821 11662 4861 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 12482 4780 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 12400 4780 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 12318 4780 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 12236 4780 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 12154 4780 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 12072 4780 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 11990 4780 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 11908 4780 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 11826 4780 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 11744 4780 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4740 11662 4780 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 12482 4699 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 12400 4699 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 12318 4699 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 12236 4699 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 12154 4699 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 12072 4699 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 11990 4699 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 11908 4699 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 11826 4699 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 11744 4699 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4659 11662 4699 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 12482 4618 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 12400 4618 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 12318 4618 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 12236 4618 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 12154 4618 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 12072 4618 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 11990 4618 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 11908 4618 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 11826 4618 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 11744 4618 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4578 11662 4618 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 12482 4537 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 12400 4537 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 12318 4537 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 12236 4537 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 12154 4537 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 12072 4537 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 11990 4537 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 11908 4537 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 11826 4537 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 11744 4537 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4497 11662 4537 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 12482 4456 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 12400 4456 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 12318 4456 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 12236 4456 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 12154 4456 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 12072 4456 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 11990 4456 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 11908 4456 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 11826 4456 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 11744 4456 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4416 11662 4456 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 12482 4375 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 12400 4375 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 12318 4375 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 12236 4375 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 12154 4375 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 12072 4375 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 11990 4375 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 11908 4375 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 11826 4375 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 11744 4375 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4335 11662 4375 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 12482 4294 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 12400 4294 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 12318 4294 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 12236 4294 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 12154 4294 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 12072 4294 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 11990 4294 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 11908 4294 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 11826 4294 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 11744 4294 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4254 11662 4294 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 12482 4213 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 12400 4213 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 12318 4213 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 12236 4213 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 12154 4213 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 12072 4213 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 11990 4213 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 11908 4213 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 11826 4213 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 11744 4213 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4173 11662 4213 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 12482 4132 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 12400 4132 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 12318 4132 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 12236 4132 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 12154 4132 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 12072 4132 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 11990 4132 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 11908 4132 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 11826 4132 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 11744 4132 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4092 11662 4132 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 12482 4051 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 12400 4051 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 12318 4051 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 12236 4051 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 12154 4051 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 12072 4051 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 11990 4051 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 11908 4051 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 11826 4051 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 11744 4051 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 4011 11662 4051 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 12482 3970 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 12400 3970 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 12318 3970 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 12236 3970 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 12154 3970 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 12072 3970 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 11990 3970 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 11908 3970 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 11826 3970 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 11744 3970 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3930 11662 3970 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 12482 3889 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 12400 3889 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 12318 3889 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 12236 3889 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 12154 3889 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 12072 3889 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 11990 3889 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 11908 3889 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 11826 3889 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 11744 3889 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3849 11662 3889 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 12482 3808 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 12400 3808 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 12318 3808 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 12236 3808 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 12154 3808 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 12072 3808 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 11990 3808 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 11908 3808 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 11826 3808 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 11744 3808 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3768 11662 3808 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 12482 3727 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 12400 3727 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 12318 3727 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 12236 3727 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 12154 3727 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 12072 3727 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 11990 3727 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 11908 3727 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 11826 3727 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 11744 3727 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3687 11662 3727 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 12482 3646 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 12400 3646 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 12318 3646 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 12236 3646 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 12154 3646 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 12072 3646 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 11990 3646 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 11908 3646 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 11826 3646 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 11744 3646 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3606 11662 3646 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 12482 3565 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 12400 3565 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 12318 3565 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 12236 3565 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 12154 3565 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 12072 3565 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 11990 3565 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 11908 3565 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 11826 3565 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 11744 3565 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3525 11662 3565 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 12482 3484 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 12400 3484 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 12318 3484 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 12236 3484 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 12154 3484 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 12072 3484 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 11990 3484 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 11908 3484 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 11826 3484 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 11744 3484 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3444 11662 3484 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 12482 3403 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 12400 3403 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 12318 3403 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 12236 3403 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 12154 3403 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 12072 3403 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 11990 3403 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 11908 3403 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 11826 3403 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 11744 3403 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3363 11662 3403 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 12482 3322 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 12400 3322 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 12318 3322 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 12236 3322 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 12154 3322 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 12072 3322 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 11990 3322 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 11908 3322 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 11826 3322 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 11744 3322 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3282 11662 3322 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 12482 3241 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 12400 3241 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 12318 3241 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 12236 3241 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 12154 3241 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 12072 3241 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 11990 3241 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 11908 3241 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 11826 3241 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 11744 3241 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3201 11662 3241 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 12482 3160 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 12400 3160 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 12318 3160 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 12236 3160 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 12154 3160 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 12072 3160 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 11990 3160 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 11908 3160 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 11826 3160 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 11744 3160 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3120 11662 3160 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 12482 3079 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 12400 3079 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 12318 3079 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 12236 3079 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 12154 3079 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 12072 3079 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 11990 3079 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 11908 3079 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 11826 3079 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 11744 3079 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 3039 11662 3079 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 12482 2998 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 12400 2998 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 12318 2998 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 12236 2998 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 12154 2998 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 12072 2998 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 11990 2998 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 11908 2998 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 11826 2998 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 11744 2998 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2958 11662 2998 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 12482 2917 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 12400 2917 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 12318 2917 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 12236 2917 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 12154 2917 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 12072 2917 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 11990 2917 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 11908 2917 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 11826 2917 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 11744 2917 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2877 11662 2917 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 12482 2836 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 12400 2836 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 12318 2836 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 12236 2836 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 12154 2836 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 12072 2836 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 11990 2836 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 11908 2836 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 11826 2836 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 11744 2836 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2796 11662 2836 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 12482 2755 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 12400 2755 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 12318 2755 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 12236 2755 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 12154 2755 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 12072 2755 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 11990 2755 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 11908 2755 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 11826 2755 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 11744 2755 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2715 11662 2755 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 12482 2674 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 12400 2674 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 12318 2674 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 12236 2674 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 12154 2674 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 12072 2674 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 11990 2674 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 11908 2674 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 11826 2674 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 11744 2674 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2634 11662 2674 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 12482 2593 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 12400 2593 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 12318 2593 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 12236 2593 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 12154 2593 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 12072 2593 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 11990 2593 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 11908 2593 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 11826 2593 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 11744 2593 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2553 11662 2593 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 12482 2512 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 12400 2512 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 12318 2512 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 12236 2512 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 12154 2512 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 12072 2512 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 11990 2512 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 11908 2512 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 11826 2512 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 11744 2512 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2472 11662 2512 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 12482 2431 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 12400 2431 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 12318 2431 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 12236 2431 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 12154 2431 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 12072 2431 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 11990 2431 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 11908 2431 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 11826 2431 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 11744 2431 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2391 11662 2431 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 12482 2350 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 12400 2350 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 12318 2350 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 12236 2350 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 12154 2350 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 12072 2350 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 11990 2350 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 11908 2350 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 11826 2350 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 11744 2350 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2310 11662 2350 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 12482 2269 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 12400 2269 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 12318 2269 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 12236 2269 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 12154 2269 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 12072 2269 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 11990 2269 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 11908 2269 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 11826 2269 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 11744 2269 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2229 11662 2269 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 12482 2188 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 12400 2188 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 12318 2188 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 12236 2188 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 12154 2188 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 12072 2188 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 11990 2188 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 11908 2188 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 11826 2188 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 11744 2188 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2148 11662 2188 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 12482 2107 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 12400 2107 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 12318 2107 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 12236 2107 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 12154 2107 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 12072 2107 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 11990 2107 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 11908 2107 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 11826 2107 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 11744 2107 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 2067 11662 2107 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 12482 2026 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 12400 2026 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 12318 2026 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 12236 2026 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 12154 2026 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 12072 2026 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 11990 2026 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 11908 2026 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 11826 2026 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 11744 2026 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1986 11662 2026 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 12482 1945 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 12400 1945 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 12318 1945 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 12236 1945 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 12154 1945 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 12072 1945 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 11990 1945 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 11908 1945 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 11826 1945 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 11744 1945 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1905 11662 1945 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 12482 1864 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 12400 1864 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 12318 1864 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 12236 1864 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 12154 1864 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 12072 1864 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 11990 1864 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 11908 1864 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 11826 1864 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 11744 1864 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1824 11662 1864 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 12482 1783 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 12400 1783 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 12318 1783 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 12236 1783 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 12154 1783 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 12072 1783 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 11990 1783 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 11908 1783 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 11826 1783 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 11744 1783 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1743 11662 1783 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 12482 1702 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 12400 1702 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 12318 1702 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 12236 1702 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 12154 1702 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 12072 1702 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 11990 1702 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 11908 1702 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 11826 1702 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 11744 1702 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1662 11662 1702 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 12482 1621 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 12400 1621 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 12318 1621 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 12236 1621 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 12154 1621 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 12072 1621 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 11990 1621 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 11908 1621 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 11826 1621 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 11744 1621 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1581 11662 1621 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 12482 1540 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 12400 1540 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 12318 1540 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 12236 1540 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 12154 1540 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 12072 1540 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 11990 1540 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 11908 1540 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 11826 1540 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 11744 1540 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1500 11662 1540 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 12482 1459 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 12400 1459 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 12318 1459 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 12236 1459 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 12154 1459 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 12072 1459 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 11990 1459 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 11908 1459 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 11826 1459 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 11744 1459 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1419 11662 1459 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 12482 1378 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 12400 1378 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 12318 1378 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 12236 1378 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 12154 1378 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 12072 1378 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 11990 1378 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 11908 1378 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 11826 1378 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 11744 1378 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1338 11662 1378 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 12482 1297 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 12400 1297 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 12318 1297 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 12236 1297 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 12154 1297 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 12072 1297 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 11990 1297 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 11908 1297 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 11826 1297 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 11744 1297 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1257 11662 1297 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 12482 1216 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 12400 1216 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 12318 1216 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 12236 1216 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 12154 1216 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 12072 1216 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 11990 1216 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 11908 1216 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 11826 1216 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 11744 1216 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1176 11662 1216 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 12482 1135 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 12400 1135 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 12318 1135 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 12236 1135 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 12154 1135 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 12072 1135 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 11990 1135 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 11908 1135 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 11826 1135 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 11744 1135 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1095 11662 1135 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 12482 1054 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 12400 1054 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 12318 1054 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 12236 1054 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 12154 1054 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 12072 1054 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 11990 1054 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 11908 1054 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 11826 1054 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 11744 1054 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 1014 11662 1054 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 12482 973 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 12400 973 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 12318 973 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 12236 973 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 12154 973 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 12072 973 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 11990 973 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 11908 973 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 11826 973 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 11744 973 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 933 11662 973 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 12482 892 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 12400 892 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 12318 892 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 12236 892 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 12154 892 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 12072 892 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 11990 892 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 11908 892 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 11826 892 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 11744 892 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 852 11662 892 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 12482 811 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 12400 811 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 12318 811 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 12236 811 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 12154 811 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 12072 811 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 11990 811 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 11908 811 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 11826 811 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 11744 811 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 771 11662 811 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 12482 730 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 12400 730 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 12318 730 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 12236 730 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 12154 730 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 12072 730 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 11990 730 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 11908 730 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 11826 730 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 11744 730 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 690 11662 730 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 12482 649 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 12400 649 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 12318 649 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 12236 649 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 12154 649 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 12072 649 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 11990 649 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 11908 649 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 11826 649 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 11744 649 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 609 11662 649 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 12482 567 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 12400 567 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 12318 567 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 12236 567 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 12154 567 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 12072 567 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 11990 567 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 11908 567 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 11826 567 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 11744 567 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 527 11662 567 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 12482 485 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 12400 485 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 12318 485 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 12236 485 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 12154 485 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 12072 485 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 11990 485 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 11908 485 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 11826 485 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 11744 485 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 445 11662 485 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 12482 403 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 12400 403 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 12318 403 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 12236 403 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 12154 403 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 12072 403 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 11990 403 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 11908 403 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 11826 403 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 11744 403 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 363 11662 403 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 12482 321 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 12400 321 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 12318 321 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 12236 321 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 12154 321 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 12072 321 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 11990 321 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 11908 321 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 11826 321 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 11744 321 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 281 11662 321 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 12482 239 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 12400 239 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 12318 239 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 12236 239 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 12154 239 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 12072 239 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 11990 239 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 11908 239 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 11826 239 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 11744 239 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 199 11662 239 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 12482 157 12522 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 12400 157 12440 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 12318 157 12358 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 12236 157 12276 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 12154 157 12194 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 12072 157 12112 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 11990 157 12030 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 11908 157 11948 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 11826 157 11866 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 11744 157 11784 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel via3 s 117 11662 157 11702 1 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal4 s 14746 6377 15000 7067 1 VSWITCH
port 59 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 1 VSWITCH
port 59 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 1 VSWITCH
port 59 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string GDS_END 25436770
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 24961600
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
