/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.ref/sky130_fd_io/cdl/sky130_ef_io.cdl