/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/sonos/begin_of_life/typical.spice