/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p25.spice