magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 222 582
<< pwell >>
rect 5 13 183 203
rect 29 -17 63 13
<< pdiff >>
rect 31 305 157 505
<< ndiode >>
rect 31 39 157 177
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 17 51 167 493
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 184 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 29 -17 63 17
rect 121 -17 155 17
<< metal1 >>
rect 0 561 184 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 0 496 184 527
rect 0 17 184 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 184 17
rect 0 -48 184 -17
<< labels >>
flabel locali s 121 85 155 119 0 FreeSans 200 0 0 0 DIODE
flabel locali s 121 357 155 391 0 FreeSans 200 0 0 0 DIODE
flabel locali s 29 357 63 391 0 FreeSans 200 0 0 0 DIODE
flabel locali s 121 425 155 459 0 FreeSans 200 0 0 0 DIODE
flabel locali s 29 425 63 459 0 FreeSans 200 0 0 0 DIODE
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 DIODE
flabel locali s 121 289 155 323 0 FreeSans 200 0 0 0 DIODE
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 DIODE
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 DIODE
flabel locali s 121 153 155 187 0 FreeSans 200 0 0 0 DIODE
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 DIODE
flabel locali s 29 85 63 119 0 FreeSans 200 0 0 0 DIODE
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 diode_2
<< properties >>
string FIXED_BBOX 0 0 184 544
string GDS_END 3957934
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3954696
string path 0.000 0.000 4.600 0.000 
<< end >>
