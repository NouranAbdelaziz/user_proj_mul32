/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/openlane/custom_cells/lef/sky130_ef_io_core.lef