/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/sonos_see_p/end_of_life.spice