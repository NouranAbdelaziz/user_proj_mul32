/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8__wafer.corner.spice