/home/nouran/user_proj_mul32/dependencies/pdks/sky130A/libs.tech/ngspice/corners/tt/leak_discrete.spice