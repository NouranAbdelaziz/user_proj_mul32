magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal4 >>
tri 1934 33739 2266 34071 se
rect 2266 34047 12734 34071
tri 12734 34047 12758 34071 sw
rect 2266 33811 2269 34047
rect 2505 33811 2589 34047
rect 2825 33811 2909 34047
rect 3145 33811 3229 34047
rect 3465 33811 3549 34047
rect 3785 33811 3869 34047
rect 4105 33811 4189 34047
rect 4425 33811 4509 34047
rect 4745 33811 4829 34047
rect 5065 33811 5149 34047
rect 5385 33811 5469 34047
rect 5705 33811 5789 34047
rect 6025 33811 6109 34047
rect 6345 33811 6429 34047
rect 6665 33811 6749 34047
rect 6985 33811 7069 34047
rect 7305 33811 7389 34047
rect 7625 33811 7709 34047
rect 7945 33811 8029 34047
rect 8265 33811 8349 34047
rect 8585 33811 8669 34047
rect 8905 33811 8989 34047
rect 9225 33811 9309 34047
rect 9545 33811 9629 34047
rect 9865 33811 9949 34047
rect 10185 33811 10269 34047
rect 10505 33811 10589 34047
rect 10825 33811 10909 34047
rect 11145 33811 11229 34047
rect 11465 33811 11549 34047
rect 11785 33811 11869 34047
rect 12105 33811 12189 34047
rect 12425 33811 12509 34047
rect 12745 33811 12758 34047
rect 2266 33739 12758 33811
tri 1726 33531 1934 33739 se
rect 1934 33531 1947 33739
tri 1614 33419 1726 33531 se
rect 1726 33503 1947 33531
rect 2183 33685 12758 33739
tri 12758 33685 13120 34047 sw
rect 2183 33531 12871 33685
rect 2183 33503 2462 33531
tri 2462 33503 2490 33531 nw
rect 1726 33419 2378 33503
tri 2378 33419 2462 33503 nw
tri 1500 33305 1614 33419 se
rect 1614 33305 1627 33419
tri 1294 33099 1500 33305 se
rect 1500 33183 1627 33305
rect 1863 33183 2142 33419
tri 2142 33183 2378 33419 nw
tri 12510 33305 12736 33531 ne
rect 12736 33449 12871 33531
rect 13107 33531 13120 33685
tri 13120 33531 13274 33685 sw
rect 13107 33449 13274 33531
rect 12736 33365 13274 33449
tri 13274 33365 13440 33531 sw
rect 12736 33305 13191 33365
rect 1500 33099 1726 33183
tri 971 32776 1294 33099 se
rect 1294 32863 1307 33099
rect 1543 32863 1726 33099
rect 1294 32776 1726 32863
tri 962 32767 971 32776 se
rect 971 32767 984 32776
tri 960 32765 962 32767 se
rect 962 32765 984 32767
rect 960 32540 984 32765
rect 1220 32767 1726 32776
tri 1726 32767 2142 33183 nw
tri 12736 33129 12912 33305 ne
rect 12912 33129 13191 33305
rect 13427 33305 13440 33365
tri 13440 33305 13500 33365 sw
rect 13427 33129 13500 33305
tri 12912 32767 13274 33129 ne
rect 13274 33045 13500 33129
tri 13500 33045 13760 33305 sw
rect 13274 32809 13511 33045
rect 13747 32809 13760 33045
rect 13274 32767 13760 32809
rect 1220 32540 1500 32767
tri 1500 32541 1726 32767 nw
tri 13274 32541 13500 32767 ne
rect 13500 32765 13760 32767
tri 13760 32765 14040 33045 sw
rect 13500 32682 14040 32765
rect 960 32456 1500 32540
rect 960 32220 984 32456
rect 1220 32220 1500 32456
rect 960 32136 1500 32220
rect 960 31900 984 32136
rect 1220 31900 1500 32136
rect 960 31816 1500 31900
rect 960 31580 984 31816
rect 1220 31580 1500 31816
rect 960 31496 1500 31580
rect 960 31260 984 31496
rect 1220 31260 1500 31496
rect 960 31176 1500 31260
rect 960 30940 984 31176
rect 1220 30940 1500 31176
rect 960 30856 1500 30940
rect 960 30620 984 30856
rect 1220 30620 1500 30856
rect 960 30536 1500 30620
rect 960 30300 984 30536
rect 1220 30300 1500 30536
rect 960 30216 1500 30300
rect 960 29980 984 30216
rect 1220 29980 1500 30216
rect 960 29896 1500 29980
rect 960 29660 984 29896
rect 1220 29660 1500 29896
rect 960 29576 1500 29660
rect 960 29340 984 29576
rect 1220 29340 1500 29576
rect 960 29256 1500 29340
rect 960 29020 984 29256
rect 1220 29020 1500 29256
rect 960 28936 1500 29020
rect 960 28700 984 28936
rect 1220 28700 1500 28936
rect 960 28616 1500 28700
rect 960 28380 984 28616
rect 1220 28380 1500 28616
rect 960 28296 1500 28380
rect 960 28060 984 28296
rect 1220 28060 1500 28296
rect 960 27976 1500 28060
rect 960 27740 984 27976
rect 1220 27740 1500 27976
rect 960 27656 1500 27740
rect 960 27420 984 27656
rect 1220 27420 1500 27656
rect 960 27336 1500 27420
rect 960 27100 984 27336
rect 1220 27100 1500 27336
rect 960 27016 1500 27100
rect 960 26780 984 27016
rect 1220 26780 1500 27016
rect 960 26696 1500 26780
rect 960 26460 984 26696
rect 1220 26460 1500 26696
rect 960 26376 1500 26460
rect 960 26140 984 26376
rect 1220 26140 1500 26376
rect 960 26056 1500 26140
rect 960 25820 984 26056
rect 1220 25820 1500 26056
rect 960 25736 1500 25820
rect 960 25500 984 25736
rect 1220 25500 1500 25736
rect 960 25416 1500 25500
rect 960 25180 984 25416
rect 1220 25180 1500 25416
rect 960 25096 1500 25180
rect 960 24860 984 25096
rect 1220 24860 1500 25096
rect 960 24776 1500 24860
rect 960 24540 984 24776
rect 1220 24540 1500 24776
rect 960 24456 1500 24540
rect 960 24220 984 24456
rect 1220 24220 1500 24456
rect 960 24136 1500 24220
rect 960 23900 984 24136
rect 1220 23900 1500 24136
rect 960 23816 1500 23900
rect 960 23580 984 23816
rect 1220 23580 1500 23816
rect 960 23496 1500 23580
rect 960 23260 984 23496
rect 1220 23260 1500 23496
rect 960 23176 1500 23260
rect 960 22940 984 23176
rect 1220 22940 1500 23176
rect 960 22856 1500 22940
rect 960 22620 984 22856
rect 1220 22620 1500 22856
rect 960 22536 1500 22620
rect 960 22300 984 22536
rect 1220 22300 1500 22536
rect 960 22216 1500 22300
rect 960 21980 984 22216
rect 1220 21980 1500 22216
rect 960 21896 1500 21980
rect 960 21660 984 21896
rect 1220 21660 1500 21896
rect 960 21576 1500 21660
rect 960 21340 984 21576
rect 1220 21340 1500 21576
rect 960 21256 1500 21340
rect 960 21020 984 21256
rect 1220 21020 1500 21256
rect 960 20936 1500 21020
rect 960 20700 984 20936
rect 1220 20700 1500 20936
rect 960 20616 1500 20700
rect 960 20380 984 20616
rect 1220 20380 1500 20616
rect 13500 32446 13780 32682
rect 14016 32446 14040 32682
rect 13500 32362 14040 32446
rect 13500 32126 13780 32362
rect 14016 32126 14040 32362
rect 13500 32042 14040 32126
rect 13500 31806 13780 32042
rect 14016 31806 14040 32042
rect 13500 31722 14040 31806
rect 13500 31486 13780 31722
rect 14016 31486 14040 31722
rect 13500 31402 14040 31486
rect 13500 31166 13780 31402
rect 14016 31166 14040 31402
rect 13500 31082 14040 31166
rect 13500 30846 13780 31082
rect 14016 30846 14040 31082
rect 13500 30762 14040 30846
rect 13500 30526 13780 30762
rect 14016 30526 14040 30762
rect 13500 30442 14040 30526
rect 13500 30206 13780 30442
rect 14016 30206 14040 30442
rect 13500 30122 14040 30206
rect 13500 29886 13780 30122
rect 14016 29886 14040 30122
rect 13500 29802 14040 29886
rect 13500 29566 13780 29802
rect 14016 29566 14040 29802
rect 13500 29482 14040 29566
rect 13500 29246 13780 29482
rect 14016 29246 14040 29482
rect 13500 29162 14040 29246
rect 13500 28926 13780 29162
rect 14016 28926 14040 29162
rect 13500 28842 14040 28926
rect 13500 28606 13780 28842
rect 14016 28606 14040 28842
rect 13500 28522 14040 28606
rect 13500 28286 13780 28522
rect 14016 28286 14040 28522
rect 13500 28202 14040 28286
rect 13500 27966 13780 28202
rect 14016 27966 14040 28202
rect 13500 27882 14040 27966
rect 13500 27646 13780 27882
rect 14016 27646 14040 27882
rect 13500 27562 14040 27646
rect 13500 27326 13780 27562
rect 14016 27326 14040 27562
rect 13500 27242 14040 27326
rect 13500 27006 13780 27242
rect 14016 27006 14040 27242
rect 13500 26922 14040 27006
rect 13500 26686 13780 26922
rect 14016 26686 14040 26922
rect 13500 26602 14040 26686
rect 13500 26366 13780 26602
rect 14016 26366 14040 26602
rect 13500 26282 14040 26366
rect 13500 26046 13780 26282
rect 14016 26046 14040 26282
rect 13500 25962 14040 26046
rect 13500 25726 13780 25962
rect 14016 25726 14040 25962
rect 13500 25642 14040 25726
rect 13500 25406 13780 25642
rect 14016 25406 14040 25642
rect 13500 25322 14040 25406
rect 13500 25086 13780 25322
rect 14016 25086 14040 25322
rect 13500 25002 14040 25086
rect 13500 24766 13780 25002
rect 14016 24766 14040 25002
rect 13500 24682 14040 24766
rect 13500 24446 13780 24682
rect 14016 24446 14040 24682
rect 13500 24362 14040 24446
rect 13500 24126 13780 24362
rect 14016 24126 14040 24362
rect 13500 24042 14040 24126
rect 13500 23806 13780 24042
rect 14016 23806 14040 24042
rect 13500 23722 14040 23806
rect 13500 23486 13780 23722
rect 14016 23486 14040 23722
rect 13500 23402 14040 23486
rect 13500 23166 13780 23402
rect 14016 23166 14040 23402
rect 13500 23082 14040 23166
rect 13500 22846 13780 23082
rect 14016 22846 14040 23082
rect 13500 22762 14040 22846
rect 13500 22526 13780 22762
rect 14016 22526 14040 22762
rect 13500 22442 14040 22526
rect 13500 22206 13780 22442
rect 14016 22206 14040 22442
rect 13500 22122 14040 22206
rect 13500 21886 13780 22122
rect 14016 21886 14040 22122
rect 13500 21802 14040 21886
rect 13500 21566 13780 21802
rect 14016 21566 14040 21802
rect 13500 21482 14040 21566
rect 13500 21246 13780 21482
rect 14016 21246 14040 21482
rect 13500 21162 14040 21246
rect 13500 20926 13780 21162
rect 14016 20926 14040 21162
rect 13500 20842 14040 20926
rect 13500 20606 13780 20842
rect 14016 20606 14040 20842
rect 13500 20522 14040 20606
rect 960 20297 1500 20380
tri 1500 20297 1724 20521 sw
tri 13276 20297 13500 20521 se
rect 13500 20297 13780 20522
tri 960 20253 1004 20297 ne
rect 1004 20295 1724 20297
tri 1724 20295 1726 20297 sw
tri 13274 20295 13276 20297 se
rect 13276 20295 13780 20297
rect 1004 20253 1726 20295
tri 1004 20017 1240 20253 ne
rect 1240 20017 1253 20253
rect 1489 20017 1726 20253
tri 1240 19757 1500 20017 ne
rect 1500 19933 1726 20017
tri 1726 19933 2088 20295 sw
rect 1500 19757 1573 19933
tri 1500 19697 1560 19757 ne
rect 1560 19697 1573 19757
rect 1809 19757 2088 19933
tri 2088 19757 2264 19933 sw
tri 12858 19879 13274 20295 se
rect 13274 20286 13780 20295
rect 14016 20297 14040 20522
rect 14016 20295 14038 20297
tri 14038 20295 14040 20297 nw
rect 14016 20286 14029 20295
tri 14029 20286 14038 20295 nw
rect 13274 20199 13942 20286
tri 13942 20199 14029 20286 nw
rect 13274 19963 13457 20199
rect 13693 19963 13706 20199
tri 13706 19963 13942 20199 nw
rect 13274 19879 13500 19963
tri 12736 19757 12858 19879 se
rect 12858 19757 13137 19879
rect 1809 19697 2264 19757
tri 1560 19531 1726 19697 ne
rect 1726 19613 2264 19697
rect 1726 19531 1893 19613
tri 1726 19377 1880 19531 ne
rect 1880 19377 1893 19531
rect 2129 19531 2264 19613
tri 2264 19531 2490 19757 sw
tri 12510 19531 12736 19757 se
rect 12736 19643 13137 19757
rect 13373 19757 13500 19879
tri 13500 19757 13706 19963 nw
rect 13373 19643 13386 19757
tri 13386 19643 13500 19757 nw
rect 12736 19559 13274 19643
rect 12736 19531 12817 19559
rect 2129 19377 12817 19531
tri 1880 19251 2006 19377 ne
rect 2006 19323 12817 19377
rect 13053 19531 13274 19559
tri 13274 19531 13386 19643 nw
rect 13053 19323 13066 19531
tri 13066 19323 13274 19531 nw
rect 2006 19251 12734 19323
tri 2006 19015 2242 19251 ne
rect 2242 19015 2255 19251
rect 2491 19015 2575 19251
rect 2811 19015 2895 19251
rect 3131 19015 3215 19251
rect 3451 19015 3535 19251
rect 3771 19015 3855 19251
rect 4091 19015 4175 19251
rect 4411 19015 4495 19251
rect 4731 19015 4815 19251
rect 5051 19015 5135 19251
rect 5371 19015 5455 19251
rect 5691 19015 5775 19251
rect 6011 19015 6095 19251
rect 6331 19015 6415 19251
rect 6651 19015 6735 19251
rect 6971 19015 7055 19251
rect 7291 19015 7375 19251
rect 7611 19015 7695 19251
rect 7931 19015 8015 19251
rect 8251 19015 8335 19251
rect 8571 19015 8655 19251
rect 8891 19015 8975 19251
rect 9211 19015 9295 19251
rect 9531 19015 9615 19251
rect 9851 19015 9935 19251
rect 10171 19015 10255 19251
rect 10491 19015 10575 19251
rect 10811 19015 10895 19251
rect 11131 19015 11215 19251
rect 11451 19015 11535 19251
rect 11771 19015 11855 19251
rect 12091 19015 12175 19251
rect 12411 19015 12495 19251
rect 12731 19015 12734 19251
tri 2242 18991 2266 19015 ne
rect 2266 18991 12734 19015
tri 12734 18991 13066 19323 nw
<< via4 >>
rect 2269 33811 2505 34047
rect 2589 33811 2825 34047
rect 2909 33811 3145 34047
rect 3229 33811 3465 34047
rect 3549 33811 3785 34047
rect 3869 33811 4105 34047
rect 4189 33811 4425 34047
rect 4509 33811 4745 34047
rect 4829 33811 5065 34047
rect 5149 33811 5385 34047
rect 5469 33811 5705 34047
rect 5789 33811 6025 34047
rect 6109 33811 6345 34047
rect 6429 33811 6665 34047
rect 6749 33811 6985 34047
rect 7069 33811 7305 34047
rect 7389 33811 7625 34047
rect 7709 33811 7945 34047
rect 8029 33811 8265 34047
rect 8349 33811 8585 34047
rect 8669 33811 8905 34047
rect 8989 33811 9225 34047
rect 9309 33811 9545 34047
rect 9629 33811 9865 34047
rect 9949 33811 10185 34047
rect 10269 33811 10505 34047
rect 10589 33811 10825 34047
rect 10909 33811 11145 34047
rect 11229 33811 11465 34047
rect 11549 33811 11785 34047
rect 11869 33811 12105 34047
rect 12189 33811 12425 34047
rect 12509 33811 12745 34047
rect 1947 33503 2183 33739
rect 1627 33183 1863 33419
rect 12871 33449 13107 33685
rect 1307 32863 1543 33099
rect 984 32540 1220 32776
rect 13191 33129 13427 33365
rect 13511 32809 13747 33045
rect 984 32220 1220 32456
rect 984 31900 1220 32136
rect 984 31580 1220 31816
rect 984 31260 1220 31496
rect 984 30940 1220 31176
rect 984 30620 1220 30856
rect 984 30300 1220 30536
rect 984 29980 1220 30216
rect 984 29660 1220 29896
rect 984 29340 1220 29576
rect 984 29020 1220 29256
rect 984 28700 1220 28936
rect 984 28380 1220 28616
rect 984 28060 1220 28296
rect 984 27740 1220 27976
rect 984 27420 1220 27656
rect 984 27100 1220 27336
rect 984 26780 1220 27016
rect 984 26460 1220 26696
rect 984 26140 1220 26376
rect 984 25820 1220 26056
rect 984 25500 1220 25736
rect 984 25180 1220 25416
rect 984 24860 1220 25096
rect 984 24540 1220 24776
rect 984 24220 1220 24456
rect 984 23900 1220 24136
rect 984 23580 1220 23816
rect 984 23260 1220 23496
rect 984 22940 1220 23176
rect 984 22620 1220 22856
rect 984 22300 1220 22536
rect 984 21980 1220 22216
rect 984 21660 1220 21896
rect 984 21340 1220 21576
rect 984 21020 1220 21256
rect 984 20700 1220 20936
rect 984 20380 1220 20616
rect 13780 32446 14016 32682
rect 13780 32126 14016 32362
rect 13780 31806 14016 32042
rect 13780 31486 14016 31722
rect 13780 31166 14016 31402
rect 13780 30846 14016 31082
rect 13780 30526 14016 30762
rect 13780 30206 14016 30442
rect 13780 29886 14016 30122
rect 13780 29566 14016 29802
rect 13780 29246 14016 29482
rect 13780 28926 14016 29162
rect 13780 28606 14016 28842
rect 13780 28286 14016 28522
rect 13780 27966 14016 28202
rect 13780 27646 14016 27882
rect 13780 27326 14016 27562
rect 13780 27006 14016 27242
rect 13780 26686 14016 26922
rect 13780 26366 14016 26602
rect 13780 26046 14016 26282
rect 13780 25726 14016 25962
rect 13780 25406 14016 25642
rect 13780 25086 14016 25322
rect 13780 24766 14016 25002
rect 13780 24446 14016 24682
rect 13780 24126 14016 24362
rect 13780 23806 14016 24042
rect 13780 23486 14016 23722
rect 13780 23166 14016 23402
rect 13780 22846 14016 23082
rect 13780 22526 14016 22762
rect 13780 22206 14016 22442
rect 13780 21886 14016 22122
rect 13780 21566 14016 21802
rect 13780 21246 14016 21482
rect 13780 20926 14016 21162
rect 13780 20606 14016 20842
rect 1253 20017 1489 20253
rect 1573 19697 1809 19933
rect 13780 20286 14016 20522
rect 13457 19963 13693 20199
rect 1893 19377 2129 19613
rect 13137 19643 13373 19879
rect 12817 19323 13053 19559
rect 2255 19015 2491 19251
rect 2575 19015 2811 19251
rect 2895 19015 3131 19251
rect 3215 19015 3451 19251
rect 3535 19015 3771 19251
rect 3855 19015 4091 19251
rect 4175 19015 4411 19251
rect 4495 19015 4731 19251
rect 4815 19015 5051 19251
rect 5135 19015 5371 19251
rect 5455 19015 5691 19251
rect 5775 19015 6011 19251
rect 6095 19015 6331 19251
rect 6415 19015 6651 19251
rect 6735 19015 6971 19251
rect 7055 19015 7291 19251
rect 7375 19015 7611 19251
rect 7695 19015 7931 19251
rect 8015 19015 8251 19251
rect 8335 19015 8571 19251
rect 8655 19015 8891 19251
rect 8975 19015 9211 19251
rect 9295 19015 9531 19251
rect 9615 19015 9851 19251
rect 9935 19015 10171 19251
rect 10255 19015 10491 19251
rect 10575 19015 10811 19251
rect 10895 19015 11131 19251
rect 11215 19015 11451 19251
rect 11535 19015 11771 19251
rect 11855 19015 12091 19251
rect 12175 19015 12411 19251
rect 12495 19015 12731 19251
<< metal5 >>
tri 1934 33739 2266 34071 se
rect 2266 34047 12734 34071
tri 12734 34047 12758 34071 sw
rect 2266 33811 2269 34047
rect 2505 33811 2589 34047
rect 2825 33811 2909 34047
rect 3145 33811 3229 34047
rect 3465 33811 3549 34047
rect 3785 33811 3869 34047
rect 4105 33811 4189 34047
rect 4425 33811 4509 34047
rect 4745 33811 4829 34047
rect 5065 33811 5149 34047
rect 5385 33811 5469 34047
rect 5705 33811 5789 34047
rect 6025 33811 6109 34047
rect 6345 33811 6429 34047
rect 6665 33811 6749 34047
rect 6985 33811 7069 34047
rect 7305 33811 7389 34047
rect 7625 33811 7709 34047
rect 7945 33811 8029 34047
rect 8265 33811 8349 34047
rect 8585 33811 8669 34047
rect 8905 33811 8989 34047
rect 9225 33811 9309 34047
rect 9545 33811 9629 34047
rect 9865 33811 9949 34047
rect 10185 33811 10269 34047
rect 10505 33811 10589 34047
rect 10825 33811 10909 34047
rect 11145 33811 11229 34047
rect 11465 33811 11549 34047
rect 11785 33811 11869 34047
rect 12105 33811 12189 34047
rect 12425 33811 12509 34047
rect 12745 33811 12758 34047
rect 2266 33739 12758 33811
tri 1731 33536 1934 33739 se
rect 1934 33536 1947 33739
tri 1614 33419 1731 33536 se
rect 1731 33503 1947 33536
rect 2183 33685 12758 33739
tri 12758 33685 13120 34047 sw
rect 2183 33683 12871 33685
rect 2183 33663 2405 33683
tri 2405 33663 2425 33683 nw
tri 12578 33663 12598 33683 ne
rect 12598 33663 12871 33683
rect 2183 33648 2390 33663
tri 2390 33648 2405 33663 nw
tri 2418 33648 2433 33663 se
rect 2433 33648 12570 33663
tri 12570 33648 12585 33663 sw
tri 12598 33648 12613 33663 ne
rect 12613 33648 12871 33663
rect 2183 33620 2362 33648
tri 2362 33620 2390 33648 nw
tri 2405 33635 2418 33648 se
rect 2418 33635 12585 33648
tri 12585 33635 12598 33648 sw
tri 12613 33635 12626 33648 ne
rect 12626 33635 12871 33648
tri 2390 33620 2405 33635 se
rect 2405 33620 12598 33635
tri 12598 33620 12613 33635 sw
tri 12626 33620 12641 33635 ne
rect 12641 33620 12871 33635
rect 2183 33592 2334 33620
tri 2334 33592 2362 33620 nw
tri 2377 33607 2390 33620 se
rect 2390 33607 12613 33620
tri 12613 33607 12626 33620 sw
tri 12641 33607 12654 33620 ne
rect 12654 33607 12871 33620
tri 2362 33592 2377 33607 se
rect 2377 33592 12626 33607
tri 12626 33592 12641 33607 sw
tri 12654 33592 12669 33607 ne
rect 12669 33592 12871 33607
rect 2183 33564 2306 33592
tri 2306 33564 2334 33592 nw
tri 2349 33579 2362 33592 se
rect 2362 33579 12641 33592
tri 12641 33579 12654 33592 sw
tri 12669 33579 12682 33592 ne
rect 12682 33579 12871 33592
tri 2334 33564 2349 33579 se
rect 2349 33564 12654 33579
tri 12654 33564 12669 33579 sw
tri 12682 33564 12697 33579 ne
rect 12697 33564 12871 33579
rect 2183 33536 2278 33564
tri 2278 33536 2306 33564 nw
tri 2321 33551 2334 33564 se
rect 2334 33551 12669 33564
tri 12669 33551 12682 33564 sw
tri 12697 33551 12710 33564 ne
rect 12710 33551 12871 33564
tri 2306 33536 2321 33551 se
rect 2321 33536 12682 33551
tri 12682 33536 12697 33551 sw
tri 12710 33536 12725 33551 ne
rect 12725 33536 12871 33551
rect 2183 33508 2250 33536
tri 2250 33508 2278 33536 nw
tri 2293 33523 2306 33536 se
rect 2306 33523 12697 33536
tri 12697 33523 12710 33536 sw
tri 12725 33523 12738 33536 ne
rect 12738 33523 12871 33536
tri 2278 33508 2293 33523 se
rect 2293 33508 12710 33523
tri 12710 33508 12725 33523 sw
tri 12738 33508 12753 33523 ne
rect 12753 33508 12871 33523
rect 2183 33503 2222 33508
rect 1731 33480 2222 33503
tri 2222 33480 2250 33508 nw
tri 2265 33495 2278 33508 se
rect 2278 33495 12725 33508
tri 12725 33495 12738 33508 sw
tri 12753 33495 12766 33508 ne
rect 12766 33495 12871 33508
tri 2250 33480 2265 33495 se
rect 2265 33480 12738 33495
tri 12738 33480 12753 33495 sw
tri 12766 33480 12781 33495 ne
rect 12781 33480 12871 33495
rect 1731 33452 2194 33480
tri 2194 33452 2222 33480 nw
tri 2237 33467 2250 33480 se
rect 2250 33467 12753 33480
tri 12753 33467 12766 33480 sw
tri 12781 33467 12794 33480 ne
rect 12794 33467 12871 33480
tri 2222 33452 2237 33467 se
rect 2237 33452 12766 33467
tri 12766 33452 12781 33467 sw
tri 12794 33452 12809 33467 ne
rect 12809 33452 12871 33467
rect 1731 33424 2166 33452
tri 2166 33424 2194 33452 nw
tri 2209 33439 2222 33452 se
rect 2222 33439 12781 33452
tri 12781 33439 12794 33452 sw
tri 12809 33439 12822 33452 ne
rect 12822 33449 12871 33452
rect 13107 33551 13120 33685
tri 13120 33551 13254 33685 sw
rect 13107 33449 13254 33551
rect 12822 33439 13254 33449
tri 2194 33424 2209 33439 se
rect 2209 33424 12794 33439
tri 12794 33424 12809 33439 sw
tri 12822 33424 12837 33439 ne
rect 12837 33424 13254 33439
rect 1731 33419 2138 33424
tri 1294 33099 1614 33419 se
rect 1614 33183 1627 33419
rect 1863 33396 2138 33419
tri 2138 33396 2166 33424 nw
tri 2181 33411 2194 33424 se
rect 2194 33411 12809 33424
tri 12809 33411 12822 33424 sw
tri 12837 33411 12850 33424 ne
rect 12850 33411 13254 33424
tri 2166 33396 2181 33411 se
rect 2181 33396 12822 33411
tri 12822 33396 12837 33411 sw
tri 12850 33396 12865 33411 ne
rect 12865 33396 13254 33411
rect 1863 33368 2110 33396
tri 2110 33368 2138 33396 nw
tri 2153 33383 2166 33396 se
rect 2166 33383 12837 33396
tri 12837 33383 12850 33396 sw
tri 12865 33383 12878 33396 ne
rect 12878 33383 13254 33396
tri 2138 33368 2153 33383 se
rect 2153 33368 12850 33383
tri 12850 33368 12865 33383 sw
tri 12878 33368 12893 33383 ne
rect 12893 33368 13254 33383
rect 1863 33340 2082 33368
tri 2082 33340 2110 33368 nw
tri 2125 33355 2138 33368 se
rect 2138 33355 12865 33368
tri 12865 33355 12878 33368 sw
tri 12893 33355 12906 33368 ne
rect 12906 33365 13254 33368
tri 13254 33365 13440 33551 sw
rect 12906 33355 13191 33365
tri 2110 33340 2125 33355 se
rect 2125 33340 12878 33355
tri 12878 33340 12893 33355 sw
tri 12906 33340 12921 33355 ne
rect 12921 33340 13191 33355
rect 1863 33312 2054 33340
tri 2054 33312 2082 33340 nw
tri 2097 33327 2110 33340 se
rect 2110 33327 12893 33340
tri 12893 33327 12906 33340 sw
tri 12921 33327 12934 33340 ne
rect 12934 33327 13191 33340
tri 2082 33312 2097 33327 se
rect 2097 33312 12906 33327
tri 12906 33312 12921 33327 sw
tri 12934 33312 12949 33327 ne
rect 12949 33312 13191 33327
rect 1863 33284 2026 33312
tri 2026 33284 2054 33312 nw
tri 2069 33299 2082 33312 se
rect 2082 33299 12921 33312
tri 12921 33299 12934 33312 sw
tri 12949 33299 12962 33312 ne
rect 12962 33299 13191 33312
tri 2054 33284 2069 33299 se
rect 2069 33284 12934 33299
tri 12934 33284 12949 33299 sw
tri 12962 33284 12977 33299 ne
rect 12977 33284 13191 33299
rect 1863 33256 1998 33284
tri 1998 33256 2026 33284 nw
tri 2041 33271 2054 33284 se
rect 2054 33271 12949 33284
tri 12949 33271 12962 33284 sw
tri 12977 33271 12990 33284 ne
rect 12990 33271 13191 33284
tri 2026 33256 2041 33271 se
rect 2041 33256 12962 33271
tri 12962 33256 12977 33271 sw
tri 12990 33256 13005 33271 ne
rect 13005 33256 13191 33271
rect 1863 33228 1970 33256
tri 1970 33228 1998 33256 nw
tri 2013 33243 2026 33256 se
rect 2026 33243 12977 33256
tri 12977 33243 12990 33256 sw
tri 13005 33243 13018 33256 ne
rect 13018 33243 13191 33256
tri 1998 33228 2013 33243 se
rect 2013 33228 12990 33243
tri 12990 33228 13005 33243 sw
tri 13018 33228 13033 33243 ne
rect 13033 33228 13191 33243
rect 1863 33200 1942 33228
tri 1942 33200 1970 33228 nw
tri 1985 33215 1998 33228 se
rect 1998 33215 13005 33228
tri 13005 33215 13018 33228 sw
tri 13033 33215 13046 33228 ne
rect 13046 33215 13191 33228
tri 1970 33200 1985 33215 se
rect 1985 33200 13018 33215
tri 13018 33200 13033 33215 sw
tri 13046 33200 13061 33215 ne
rect 13061 33200 13191 33215
rect 1863 33183 1914 33200
rect 1614 33172 1914 33183
tri 1914 33172 1942 33200 nw
tri 1957 33187 1970 33200 se
rect 1970 33187 13033 33200
tri 13033 33187 13046 33200 sw
tri 13061 33187 13074 33200 ne
rect 13074 33187 13191 33200
tri 1942 33172 1957 33187 se
rect 1957 33172 13046 33187
tri 13046 33172 13061 33187 sw
tri 13074 33172 13089 33187 ne
rect 13089 33172 13191 33187
rect 1614 33144 1886 33172
tri 1886 33144 1914 33172 nw
tri 1929 33159 1942 33172 se
rect 1942 33159 13061 33172
tri 13061 33159 13074 33172 sw
tri 13089 33159 13102 33172 ne
rect 13102 33159 13191 33172
tri 1914 33144 1929 33159 se
rect 1929 33144 13074 33159
tri 13074 33144 13089 33159 sw
tri 13102 33144 13117 33159 ne
rect 13117 33144 13191 33159
rect 1614 33116 1858 33144
tri 1858 33116 1886 33144 nw
tri 1901 33131 1914 33144 se
rect 1914 33131 13089 33144
tri 13089 33131 13102 33144 sw
tri 13117 33131 13130 33144 ne
rect 13130 33131 13191 33144
tri 1886 33116 1901 33131 se
rect 1901 33116 13102 33131
tri 13102 33116 13117 33131 sw
tri 13130 33116 13145 33131 ne
rect 13145 33129 13191 33131
rect 13427 33129 13440 33365
rect 13145 33116 13440 33129
rect 1614 33099 1830 33116
tri 1199 33004 1294 33099 se
rect 1294 33004 1307 33099
tri 971 32776 1199 33004 se
rect 1199 32863 1307 33004
rect 1543 33088 1830 33099
tri 1830 33088 1858 33116 nw
tri 1873 33103 1886 33116 se
rect 1886 33103 13117 33116
tri 13117 33103 13130 33116 sw
tri 13145 33103 13158 33116 ne
rect 13158 33103 13440 33116
tri 1858 33088 1873 33103 se
rect 1873 33088 13130 33103
tri 13130 33088 13145 33103 sw
tri 13158 33088 13173 33103 ne
rect 13173 33088 13440 33103
rect 1543 33060 1802 33088
tri 1802 33060 1830 33088 nw
tri 1845 33075 1858 33088 se
rect 1858 33075 13145 33088
tri 13145 33075 13158 33088 sw
tri 13173 33075 13186 33088 ne
rect 13186 33075 13440 33088
tri 1830 33060 1845 33075 se
rect 1845 33060 13158 33075
tri 13158 33060 13173 33075 sw
tri 13186 33060 13201 33075 ne
rect 13201 33060 13440 33075
rect 1543 33032 1774 33060
tri 1774 33032 1802 33060 nw
tri 1817 33047 1830 33060 se
rect 1830 33047 13173 33060
tri 13173 33047 13186 33060 sw
tri 13201 33047 13214 33060 ne
rect 13214 33047 13440 33060
tri 1802 33032 1817 33047 se
rect 1817 33032 13186 33047
tri 13186 33032 13201 33047 sw
tri 13214 33032 13229 33047 ne
rect 13229 33045 13440 33047
tri 13440 33045 13760 33365 sw
rect 13229 33032 13511 33045
rect 1543 33004 1746 33032
tri 1746 33004 1774 33032 nw
tri 1789 33019 1802 33032 se
rect 1802 33019 13201 33032
tri 13201 33019 13214 33032 sw
tri 13229 33019 13242 33032 ne
rect 13242 33019 13511 33032
tri 1774 33004 1789 33019 se
rect 1789 33004 13214 33019
tri 13214 33004 13229 33019 sw
tri 13242 33004 13257 33019 ne
rect 13257 33004 13511 33019
rect 1543 32976 1718 33004
tri 1718 32976 1746 33004 nw
tri 1761 32991 1774 33004 se
rect 1774 32991 13229 33004
tri 13229 32991 13242 33004 sw
tri 13257 32991 13270 33004 ne
rect 13270 32991 13511 33004
tri 1746 32976 1761 32991 se
rect 1761 32976 13242 32991
tri 13242 32976 13257 32991 sw
tri 13270 32976 13285 32991 ne
rect 13285 32976 13511 32991
rect 1543 32948 1690 32976
tri 1690 32948 1718 32976 nw
tri 1733 32963 1746 32976 se
rect 1746 32963 13257 32976
tri 13257 32963 13270 32976 sw
tri 13285 32963 13298 32976 ne
rect 13298 32963 13511 32976
tri 1718 32948 1733 32963 se
rect 1733 32948 13270 32963
tri 13270 32948 13285 32963 sw
tri 13298 32948 13313 32963 ne
rect 13313 32948 13511 32963
rect 1543 32920 1662 32948
tri 1662 32920 1690 32948 nw
tri 1705 32935 1718 32948 se
rect 1718 32935 13285 32948
tri 13285 32935 13298 32948 sw
tri 13313 32935 13326 32948 ne
rect 13326 32935 13511 32948
tri 1690 32920 1705 32935 se
rect 1705 32920 13298 32935
tri 13298 32920 13313 32935 sw
tri 13326 32920 13341 32935 ne
rect 13341 32920 13511 32935
rect 1543 32892 1634 32920
tri 1634 32892 1662 32920 nw
tri 1677 32907 1690 32920 se
rect 1690 32907 13313 32920
tri 13313 32907 13326 32920 sw
tri 13341 32907 13354 32920 ne
rect 13354 32907 13511 32920
tri 1662 32892 1677 32907 se
rect 1677 32892 13326 32907
tri 13326 32892 13341 32907 sw
tri 13354 32892 13369 32907 ne
rect 13369 32892 13511 32907
rect 1543 32864 1606 32892
tri 1606 32864 1634 32892 nw
tri 1649 32879 1662 32892 se
rect 1662 32879 13341 32892
tri 13341 32879 13354 32892 sw
tri 13369 32879 13382 32892 ne
rect 13382 32879 13511 32892
tri 1634 32864 1649 32879 se
rect 1649 32864 13354 32879
tri 13354 32864 13369 32879 sw
tri 13382 32864 13397 32879 ne
rect 13397 32864 13511 32879
rect 1543 32863 1578 32864
rect 1199 32836 1578 32863
tri 1578 32836 1606 32864 nw
tri 1621 32851 1634 32864 se
rect 1634 32851 13369 32864
tri 13369 32851 13382 32864 sw
tri 13397 32851 13410 32864 ne
rect 13410 32851 13511 32864
tri 1606 32836 1621 32851 se
rect 1621 32836 13382 32851
tri 13382 32836 13397 32851 sw
tri 13410 32836 13425 32851 ne
rect 13425 32836 13511 32851
rect 1199 32808 1550 32836
tri 1550 32808 1578 32836 nw
tri 1593 32823 1606 32836 se
rect 1606 32823 13397 32836
tri 13397 32823 13410 32836 sw
tri 13425 32823 13438 32836 ne
rect 13438 32823 13511 32836
tri 1578 32808 1593 32823 se
rect 1593 32808 13410 32823
tri 13410 32808 13425 32823 sw
tri 13438 32808 13453 32823 ne
rect 13453 32809 13511 32823
rect 13747 33019 13760 33045
tri 13760 33019 13786 33045 sw
rect 13747 32809 13786 33019
rect 13453 32808 13786 32809
rect 1199 32780 1522 32808
tri 1522 32780 1550 32808 nw
tri 1565 32795 1578 32808 se
rect 1578 32795 13425 32808
tri 13425 32795 13438 32808 sw
tri 13453 32795 13466 32808 ne
rect 13466 32795 13786 32808
tri 1550 32780 1565 32795 se
rect 1565 32780 13438 32795
tri 13438 32780 13453 32795 sw
tri 13466 32780 13481 32795 ne
rect 13481 32780 13786 32795
rect 1199 32776 1507 32780
tri 960 32765 971 32776 se
rect 971 32765 984 32776
rect 960 32540 984 32765
rect 1220 32765 1507 32776
tri 1507 32765 1522 32780 nw
tri 1537 32767 1550 32780 se
rect 1550 32767 13453 32780
tri 13453 32767 13466 32780 sw
tri 13481 32767 13494 32780 ne
rect 13494 32767 13786 32780
tri 1535 32765 1537 32767 se
rect 1537 32765 13466 32767
tri 13466 32765 13468 32767 sw
tri 13494 32765 13496 32767 ne
rect 13496 32765 13786 32767
tri 13786 32765 14040 33019 sw
rect 1220 32752 1494 32765
tri 1494 32752 1507 32765 nw
tri 1522 32752 1535 32765 se
rect 1535 32752 13468 32765
tri 13468 32752 13481 32765 sw
tri 13496 32752 13509 32765 ne
rect 13509 32752 14040 32765
rect 1220 32724 1466 32752
tri 1466 32724 1494 32752 nw
tri 1509 32739 1522 32752 se
rect 1522 32739 13481 32752
tri 13481 32739 13494 32752 sw
tri 13509 32739 13522 32752 ne
rect 13522 32739 14040 32752
tri 1494 32724 1509 32739 se
rect 1509 32724 13494 32739
tri 13494 32724 13509 32739 sw
tri 13522 32724 13537 32739 ne
rect 13537 32724 14040 32739
rect 1220 32696 1438 32724
tri 1438 32696 1466 32724 nw
tri 1481 32711 1494 32724 se
rect 1494 32711 13509 32724
tri 13509 32711 13522 32724 sw
tri 13537 32711 13550 32724 ne
rect 13550 32711 14040 32724
tri 1466 32696 1481 32711 se
rect 1481 32696 13522 32711
tri 13522 32696 13537 32711 sw
tri 13550 32696 13565 32711 ne
rect 13565 32696 14040 32711
rect 1220 32668 1410 32696
tri 1410 32668 1438 32696 nw
tri 1453 32683 1466 32696 se
rect 1466 32683 13537 32696
tri 13537 32683 13550 32696 sw
tri 13565 32683 13578 32696 ne
rect 13578 32683 14040 32696
tri 1438 32668 1453 32683 se
rect 1453 32668 13550 32683
tri 13550 32668 13565 32683 sw
tri 13578 32668 13593 32683 ne
rect 13593 32682 14040 32683
rect 13593 32668 13780 32682
rect 1220 32640 1382 32668
tri 1382 32640 1410 32668 nw
tri 1425 32655 1438 32668 se
rect 1438 32655 13565 32668
tri 13565 32655 13578 32668 sw
tri 13593 32657 13604 32668 ne
rect 13604 32657 13780 32668
tri 13604 32655 13606 32657 ne
rect 13606 32655 13780 32657
tri 1410 32640 1425 32655 se
rect 1425 32640 13578 32655
tri 13578 32640 13593 32655 sw
tri 13606 32640 13621 32655 ne
rect 13621 32640 13780 32655
rect 1220 32612 1354 32640
tri 1354 32612 1382 32640 nw
tri 1399 32629 1410 32640 se
rect 1410 32629 13593 32640
tri 13593 32629 13604 32640 sw
tri 13621 32637 13624 32640 ne
tri 1382 32612 1399 32629 se
rect 1399 32612 13604 32629
rect 1220 32540 1334 32612
tri 1334 32592 1354 32612 nw
tri 1362 32592 1382 32612 se
rect 1382 32592 13604 32612
rect 960 32456 1334 32540
rect 960 32220 984 32456
rect 1220 32220 1334 32456
rect 960 32136 1334 32220
rect 960 31900 984 32136
rect 1220 31900 1334 32136
rect 960 31816 1334 31900
rect 960 31580 984 31816
rect 1220 31580 1334 31816
rect 960 31496 1334 31580
rect 960 31260 984 31496
rect 1220 31260 1334 31496
rect 960 31176 1334 31260
rect 960 30940 984 31176
rect 1220 30940 1334 31176
rect 960 30856 1334 30940
rect 960 30620 984 30856
rect 1220 30620 1334 30856
rect 960 30536 1334 30620
rect 960 30300 984 30536
rect 1220 30300 1334 30536
rect 960 30216 1334 30300
rect 960 29980 984 30216
rect 1220 29980 1334 30216
rect 960 29896 1334 29980
rect 960 29660 984 29896
rect 1220 29660 1334 29896
rect 960 29576 1334 29660
rect 960 29340 984 29576
rect 1220 29340 1334 29576
rect 960 29256 1334 29340
rect 960 29020 984 29256
rect 1220 29020 1334 29256
rect 960 28936 1334 29020
rect 960 28700 984 28936
rect 1220 28700 1334 28936
rect 960 28616 1334 28700
rect 960 28380 984 28616
rect 1220 28380 1334 28616
rect 960 28296 1334 28380
rect 960 28060 984 28296
rect 1220 28060 1334 28296
rect 960 27976 1334 28060
rect 960 27740 984 27976
rect 1220 27740 1334 27976
rect 960 27656 1334 27740
rect 960 27420 984 27656
rect 1220 27420 1334 27656
rect 960 27336 1334 27420
rect 960 27100 984 27336
rect 1220 27100 1334 27336
rect 960 27016 1334 27100
rect 960 26780 984 27016
rect 1220 26780 1334 27016
rect 960 26696 1334 26780
rect 960 26460 984 26696
rect 1220 26460 1334 26696
rect 960 26376 1334 26460
rect 960 26140 984 26376
rect 1220 26140 1334 26376
rect 960 26056 1334 26140
rect 960 25820 984 26056
rect 1220 25820 1334 26056
rect 960 25736 1334 25820
rect 960 25500 984 25736
rect 1220 25500 1334 25736
rect 960 25416 1334 25500
rect 960 25180 984 25416
rect 1220 25180 1334 25416
rect 960 25096 1334 25180
rect 960 24860 984 25096
rect 1220 24860 1334 25096
rect 960 24776 1334 24860
rect 960 24540 984 24776
rect 1220 24540 1334 24776
rect 960 24456 1334 24540
rect 960 24220 984 24456
rect 1220 24220 1334 24456
rect 960 24136 1334 24220
rect 960 23900 984 24136
rect 1220 23900 1334 24136
rect 960 23816 1334 23900
rect 960 23580 984 23816
rect 1220 23580 1334 23816
rect 960 23496 1334 23580
rect 960 23260 984 23496
rect 1220 23260 1334 23496
rect 960 23176 1334 23260
rect 960 22940 984 23176
rect 1220 22940 1334 23176
rect 960 22856 1334 22940
rect 960 22620 984 22856
rect 1220 22620 1334 22856
rect 960 22536 1334 22620
rect 960 22300 984 22536
rect 1220 22300 1334 22536
rect 960 22216 1334 22300
rect 960 21980 984 22216
rect 1220 21980 1334 22216
rect 960 21896 1334 21980
rect 960 21660 984 21896
rect 1220 21660 1334 21896
rect 960 21576 1334 21660
rect 960 21340 984 21576
rect 1220 21340 1334 21576
rect 960 21256 1334 21340
rect 960 21020 984 21256
rect 1220 21020 1334 21256
rect 960 20936 1334 21020
rect 960 20700 984 20936
rect 1220 20700 1334 20936
rect 960 20616 1334 20700
rect 960 20380 984 20616
rect 1220 20503 1334 20616
tri 1354 32584 1362 32592 se
rect 1362 32584 13604 32592
rect 1354 20528 13604 32584
tri 1354 20520 1362 20528 ne
rect 1362 20520 13604 20528
tri 1334 20503 1351 20520 sw
tri 1362 20503 1379 20520 ne
rect 1379 20503 13604 20520
rect 1220 20500 1351 20503
tri 1351 20500 1354 20503 sw
tri 1379 20500 1382 20503 ne
rect 1382 20500 13604 20503
rect 1220 20475 1354 20500
tri 1354 20475 1379 20500 sw
tri 1382 20475 1407 20500 ne
rect 1407 20475 13604 20500
rect 1220 20447 1379 20475
tri 1379 20447 1407 20475 sw
tri 1407 20473 1409 20475 ne
rect 1409 20473 13604 20475
tri 1409 20447 1435 20473 ne
rect 1435 20447 13578 20473
tri 13578 20447 13604 20473 nw
rect 13624 32446 13780 32640
rect 14016 32446 14040 32682
rect 13624 32362 14040 32446
rect 13624 32126 13780 32362
rect 14016 32126 14040 32362
rect 13624 32042 14040 32126
rect 13624 31806 13780 32042
rect 14016 31806 14040 32042
rect 13624 31722 14040 31806
rect 13624 31486 13780 31722
rect 14016 31486 14040 31722
rect 13624 31402 14040 31486
rect 13624 31166 13780 31402
rect 14016 31166 14040 31402
rect 13624 31082 14040 31166
rect 13624 30846 13780 31082
rect 14016 30846 14040 31082
rect 13624 30762 14040 30846
rect 13624 30526 13780 30762
rect 14016 30526 14040 30762
rect 13624 30442 14040 30526
rect 13624 30206 13780 30442
rect 14016 30206 14040 30442
rect 13624 30122 14040 30206
rect 13624 29886 13780 30122
rect 14016 29886 14040 30122
rect 13624 29802 14040 29886
rect 13624 29566 13780 29802
rect 14016 29566 14040 29802
rect 13624 29482 14040 29566
rect 13624 29246 13780 29482
rect 14016 29246 14040 29482
rect 13624 29162 14040 29246
rect 13624 28926 13780 29162
rect 14016 28926 14040 29162
rect 13624 28842 14040 28926
rect 13624 28606 13780 28842
rect 14016 28606 14040 28842
rect 13624 28522 14040 28606
rect 13624 28286 13780 28522
rect 14016 28286 14040 28522
rect 13624 28202 14040 28286
rect 13624 27966 13780 28202
rect 14016 27966 14040 28202
rect 13624 27882 14040 27966
rect 13624 27646 13780 27882
rect 14016 27646 14040 27882
rect 13624 27562 14040 27646
rect 13624 27326 13780 27562
rect 14016 27326 14040 27562
rect 13624 27242 14040 27326
rect 13624 27006 13780 27242
rect 14016 27006 14040 27242
rect 13624 26922 14040 27006
rect 13624 26686 13780 26922
rect 14016 26686 14040 26922
rect 13624 26602 14040 26686
rect 13624 26366 13780 26602
rect 14016 26366 14040 26602
rect 13624 26282 14040 26366
rect 13624 26046 13780 26282
rect 14016 26046 14040 26282
rect 13624 25962 14040 26046
rect 13624 25726 13780 25962
rect 14016 25726 14040 25962
rect 13624 25642 14040 25726
rect 13624 25406 13780 25642
rect 14016 25406 14040 25642
rect 13624 25322 14040 25406
rect 13624 25086 13780 25322
rect 14016 25086 14040 25322
rect 13624 25002 14040 25086
rect 13624 24766 13780 25002
rect 14016 24766 14040 25002
rect 13624 24682 14040 24766
rect 13624 24446 13780 24682
rect 14016 24446 14040 24682
rect 13624 24362 14040 24446
rect 13624 24126 13780 24362
rect 14016 24126 14040 24362
rect 13624 24042 14040 24126
rect 13624 23806 13780 24042
rect 14016 23806 14040 24042
rect 13624 23722 14040 23806
rect 13624 23486 13780 23722
rect 14016 23486 14040 23722
rect 13624 23402 14040 23486
rect 13624 23166 13780 23402
rect 14016 23166 14040 23402
rect 13624 23082 14040 23166
rect 13624 22846 13780 23082
rect 14016 22846 14040 23082
rect 13624 22762 14040 22846
rect 13624 22526 13780 22762
rect 14016 22526 14040 22762
rect 13624 22442 14040 22526
rect 13624 22206 13780 22442
rect 14016 22206 14040 22442
rect 13624 22122 14040 22206
rect 13624 21886 13780 22122
rect 14016 21886 14040 22122
rect 13624 21802 14040 21886
rect 13624 21566 13780 21802
rect 14016 21566 14040 21802
rect 13624 21482 14040 21566
rect 13624 21246 13780 21482
rect 14016 21246 14040 21482
rect 13624 21162 14040 21246
rect 13624 20926 13780 21162
rect 14016 20926 14040 21162
rect 13624 20842 14040 20926
rect 13624 20606 13780 20842
rect 14016 20606 14040 20842
rect 13624 20522 14040 20606
tri 13606 20447 13624 20465 se
rect 13624 20447 13780 20522
rect 1220 20419 1407 20447
tri 1407 20419 1435 20447 sw
tri 1435 20445 1437 20447 ne
rect 1437 20445 13576 20447
tri 13576 20445 13578 20447 nw
tri 13604 20445 13606 20447 se
rect 13606 20445 13780 20447
tri 1437 20419 1463 20445 ne
rect 1463 20419 13550 20445
tri 13550 20419 13576 20445 nw
tri 13578 20419 13604 20445 se
rect 13604 20419 13780 20445
rect 1220 20391 1435 20419
tri 1435 20391 1463 20419 sw
tri 1463 20417 1465 20419 ne
rect 1465 20417 13548 20419
tri 13548 20417 13550 20419 nw
tri 13576 20417 13578 20419 se
rect 13578 20417 13780 20419
tri 1465 20391 1491 20417 ne
rect 1491 20391 13522 20417
tri 13522 20391 13548 20417 nw
tri 13550 20391 13576 20417 se
rect 13576 20391 13780 20417
rect 1220 20380 1463 20391
rect 960 20363 1463 20380
tri 1463 20363 1491 20391 sw
tri 1491 20389 1493 20391 ne
rect 1493 20389 13520 20391
tri 13520 20389 13522 20391 nw
tri 13548 20389 13550 20391 se
rect 13550 20389 13780 20391
tri 1493 20363 1519 20389 ne
rect 1519 20363 13494 20389
tri 13494 20363 13520 20389 nw
tri 13522 20363 13548 20389 se
rect 13548 20363 13780 20389
rect 960 20335 1491 20363
tri 1491 20335 1519 20363 sw
tri 1519 20361 1521 20363 ne
rect 1521 20361 13492 20363
tri 13492 20361 13494 20363 nw
tri 13520 20361 13522 20363 se
rect 13522 20361 13780 20363
tri 1521 20335 1547 20361 ne
rect 1547 20335 13466 20361
tri 13466 20335 13492 20361 nw
tri 13494 20335 13520 20361 se
rect 13520 20335 13780 20361
rect 960 20307 1519 20335
tri 1519 20307 1547 20335 sw
tri 1547 20333 1549 20335 ne
rect 1549 20333 13464 20335
tri 13464 20333 13466 20335 nw
tri 13492 20333 13494 20335 se
rect 13494 20333 13780 20335
tri 1549 20307 1575 20333 ne
rect 1575 20307 13438 20333
tri 13438 20307 13464 20333 nw
tri 13466 20307 13492 20333 se
rect 13492 20307 13780 20333
rect 960 20297 1547 20307
tri 1547 20297 1557 20307 sw
tri 1575 20305 1577 20307 ne
rect 1577 20305 13436 20307
tri 13436 20305 13438 20307 nw
tri 13464 20305 13466 20307 se
rect 13466 20305 13780 20307
tri 1577 20297 1585 20305 ne
rect 1585 20297 13428 20305
tri 13428 20297 13436 20305 nw
tri 13456 20297 13464 20305 se
rect 13464 20297 13780 20305
tri 960 20279 978 20297 ne
rect 978 20279 1557 20297
tri 1557 20279 1575 20297 sw
tri 1585 20279 1603 20297 ne
rect 1603 20279 13410 20297
tri 13410 20279 13428 20297 nw
tri 13438 20279 13456 20297 se
rect 13456 20286 13780 20297
rect 14016 20297 14040 20522
rect 14016 20286 14020 20297
rect 13456 20279 14020 20286
tri 978 20251 1006 20279 ne
rect 1006 20253 1575 20279
rect 1006 20251 1253 20253
tri 1006 20223 1034 20251 ne
rect 1034 20223 1253 20251
tri 1034 20195 1062 20223 ne
rect 1062 20195 1253 20223
tri 1062 20167 1090 20195 ne
rect 1090 20167 1253 20195
tri 1090 20139 1118 20167 ne
rect 1118 20139 1253 20167
tri 1118 20111 1146 20139 ne
rect 1146 20111 1253 20139
tri 1146 20083 1174 20111 ne
rect 1174 20083 1253 20111
tri 1174 20055 1202 20083 ne
rect 1202 20055 1253 20083
tri 1202 20027 1230 20055 ne
rect 1230 20027 1253 20055
tri 1230 20017 1240 20027 ne
rect 1240 20017 1253 20027
rect 1489 20251 1575 20253
tri 1575 20251 1603 20279 sw
tri 1603 20277 1605 20279 ne
rect 1605 20277 13408 20279
tri 13408 20277 13410 20279 nw
tri 13436 20277 13438 20279 se
rect 13438 20277 14020 20279
tri 14020 20277 14040 20297 nw
tri 1605 20251 1631 20277 ne
rect 1631 20251 13382 20277
tri 13382 20251 13408 20277 nw
tri 13410 20251 13436 20277 se
rect 13436 20251 13992 20277
rect 1489 20223 1603 20251
tri 1603 20223 1631 20251 sw
tri 1631 20249 1633 20251 ne
rect 1633 20249 13380 20251
tri 13380 20249 13382 20251 nw
tri 13408 20249 13410 20251 se
rect 13410 20249 13992 20251
tri 13992 20249 14020 20277 nw
tri 1633 20223 1659 20249 ne
rect 1659 20223 13354 20249
tri 13354 20223 13380 20249 nw
tri 13382 20223 13408 20249 se
rect 13408 20223 13964 20249
rect 1489 20195 1631 20223
tri 1631 20195 1659 20223 sw
tri 1659 20221 1661 20223 ne
rect 1661 20221 13352 20223
tri 13352 20221 13354 20223 nw
tri 13380 20221 13382 20223 se
rect 13382 20221 13964 20223
tri 13964 20221 13992 20249 nw
tri 1661 20195 1687 20221 ne
rect 1687 20195 13326 20221
tri 13326 20195 13352 20221 nw
tri 13354 20195 13380 20221 se
rect 13380 20199 13936 20221
rect 13380 20195 13457 20199
rect 1489 20167 1659 20195
tri 1659 20167 1687 20195 sw
tri 1687 20193 1689 20195 ne
rect 1689 20193 13324 20195
tri 13324 20193 13326 20195 nw
tri 13352 20193 13354 20195 se
rect 13354 20193 13457 20195
tri 1689 20167 1715 20193 ne
rect 1715 20167 13298 20193
tri 13298 20167 13324 20193 nw
tri 13326 20167 13352 20193 se
rect 13352 20167 13457 20193
rect 1489 20139 1687 20167
tri 1687 20139 1715 20167 sw
tri 1715 20165 1717 20167 ne
rect 1717 20165 13296 20167
tri 13296 20165 13298 20167 nw
tri 13324 20165 13326 20167 se
rect 13326 20165 13457 20167
tri 1717 20139 1743 20165 ne
rect 1743 20139 13270 20165
tri 13270 20139 13296 20165 nw
tri 13298 20139 13324 20165 se
rect 13324 20139 13457 20165
rect 1489 20111 1715 20139
tri 1715 20111 1743 20139 sw
tri 1743 20137 1745 20139 ne
rect 1745 20137 13268 20139
tri 13268 20137 13270 20139 nw
tri 13296 20137 13298 20139 se
rect 13298 20137 13457 20139
tri 1745 20111 1771 20137 ne
rect 1771 20111 13242 20137
tri 13242 20111 13268 20137 nw
tri 13270 20111 13296 20137 se
rect 13296 20111 13457 20137
rect 1489 20083 1743 20111
tri 1743 20083 1771 20111 sw
tri 1771 20109 1773 20111 ne
rect 1773 20109 13240 20111
tri 13240 20109 13242 20111 nw
tri 13268 20109 13270 20111 se
rect 13270 20109 13457 20111
tri 1773 20083 1799 20109 ne
rect 1799 20083 13214 20109
tri 13214 20083 13240 20109 nw
tri 13242 20083 13268 20109 se
rect 13268 20083 13457 20109
rect 1489 20055 1771 20083
tri 1771 20055 1799 20083 sw
tri 1799 20081 1801 20083 ne
rect 1801 20081 13212 20083
tri 13212 20081 13214 20083 nw
tri 13240 20081 13242 20083 se
rect 13242 20081 13457 20083
tri 1801 20055 1827 20081 ne
rect 1827 20055 13186 20081
tri 13186 20055 13212 20081 nw
tri 13214 20055 13240 20081 se
rect 13240 20055 13457 20081
rect 1489 20027 1799 20055
tri 1799 20027 1827 20055 sw
tri 1827 20053 1829 20055 ne
rect 1829 20053 13184 20055
tri 13184 20053 13186 20055 nw
tri 13212 20053 13214 20055 se
rect 13214 20053 13457 20055
tri 1829 20027 1855 20053 ne
rect 1855 20027 13158 20053
tri 13158 20027 13184 20053 nw
tri 13186 20027 13212 20053 se
rect 13212 20027 13457 20053
rect 1489 20017 1827 20027
tri 1240 19999 1258 20017 ne
rect 1258 19999 1827 20017
tri 1827 19999 1855 20027 sw
tri 1855 20025 1857 20027 ne
rect 1857 20025 13156 20027
tri 13156 20025 13158 20027 nw
tri 13184 20025 13186 20027 se
rect 13186 20025 13457 20027
tri 1857 19999 1883 20025 ne
rect 1883 19999 13130 20025
tri 13130 19999 13156 20025 nw
tri 13158 19999 13184 20025 se
rect 13184 19999 13457 20025
tri 1258 19971 1286 19999 ne
rect 1286 19971 1855 19999
tri 1855 19971 1883 19999 sw
tri 1883 19997 1885 19999 ne
rect 1885 19997 13128 19999
tri 13128 19997 13130 19999 nw
tri 13156 19997 13158 19999 se
rect 13158 19997 13457 19999
tri 1885 19971 1911 19997 ne
rect 1911 19971 13102 19997
tri 13102 19971 13128 19997 nw
tri 13130 19971 13156 19997 se
rect 13156 19971 13457 19997
tri 1286 19943 1314 19971 ne
rect 1314 19943 1883 19971
tri 1883 19943 1911 19971 sw
tri 1911 19969 1913 19971 ne
rect 1913 19969 13100 19971
tri 13100 19969 13102 19971 nw
tri 13128 19969 13130 19971 se
rect 13130 19969 13457 19971
tri 1913 19943 1939 19969 ne
rect 1939 19943 13074 19969
tri 13074 19943 13100 19969 nw
tri 13102 19943 13128 19969 se
rect 13128 19963 13457 19969
rect 13693 20193 13936 20199
tri 13936 20193 13964 20221 nw
rect 13693 20165 13908 20193
tri 13908 20165 13936 20193 nw
rect 13693 20137 13880 20165
tri 13880 20137 13908 20165 nw
rect 13693 20109 13852 20137
tri 13852 20109 13880 20137 nw
rect 13693 20081 13824 20109
tri 13824 20081 13852 20109 nw
rect 13693 20053 13796 20081
tri 13796 20053 13824 20081 nw
rect 13693 20025 13768 20053
tri 13768 20025 13796 20053 nw
rect 13693 19997 13740 20025
tri 13740 19997 13768 20025 nw
rect 13693 19969 13712 19997
tri 13712 19969 13740 19997 nw
rect 13693 19963 13706 19969
tri 13706 19963 13712 19969 nw
rect 13128 19943 13684 19963
tri 1314 19915 1342 19943 ne
rect 1342 19933 1911 19943
rect 1342 19915 1573 19933
tri 1342 19887 1370 19915 ne
rect 1370 19887 1573 19915
tri 1370 19859 1398 19887 ne
rect 1398 19859 1573 19887
tri 1398 19831 1426 19859 ne
rect 1426 19831 1573 19859
tri 1426 19803 1454 19831 ne
rect 1454 19803 1573 19831
tri 1454 19775 1482 19803 ne
rect 1482 19775 1573 19803
tri 1482 19747 1510 19775 ne
rect 1510 19747 1573 19775
tri 1510 19719 1538 19747 ne
rect 1538 19719 1573 19747
tri 1538 19691 1566 19719 ne
rect 1566 19697 1573 19719
rect 1809 19915 1911 19933
tri 1911 19915 1939 19943 sw
tri 1939 19941 1941 19943 ne
rect 1941 19941 13072 19943
tri 13072 19941 13074 19943 nw
tri 13100 19941 13102 19943 se
rect 13102 19941 13684 19943
tri 13684 19941 13706 19963 nw
tri 1941 19915 1967 19941 ne
rect 1967 19915 13046 19941
tri 13046 19915 13072 19941 nw
tri 13074 19915 13100 19941 se
rect 13100 19915 13656 19941
rect 1809 19887 1939 19915
tri 1939 19887 1967 19915 sw
tri 1967 19913 1969 19915 ne
rect 1969 19913 13044 19915
tri 13044 19913 13046 19915 nw
tri 13072 19913 13074 19915 se
rect 13074 19913 13656 19915
tri 13656 19913 13684 19941 nw
tri 1969 19887 1995 19913 ne
rect 1995 19887 13018 19913
tri 13018 19887 13044 19913 nw
tri 13046 19887 13072 19913 se
rect 13072 19887 13628 19913
rect 1809 19859 1967 19887
tri 1967 19859 1995 19887 sw
tri 1995 19885 1997 19887 ne
rect 1997 19885 13016 19887
tri 13016 19885 13018 19887 nw
tri 13044 19885 13046 19887 se
rect 13046 19885 13628 19887
tri 13628 19885 13656 19913 nw
tri 1997 19859 2023 19885 ne
rect 2023 19859 12990 19885
tri 12990 19859 13016 19885 nw
tri 13018 19859 13044 19885 se
rect 13044 19879 13600 19885
rect 13044 19859 13137 19879
rect 1809 19831 1995 19859
tri 1995 19831 2023 19859 sw
tri 2023 19857 2025 19859 ne
rect 2025 19857 12988 19859
tri 12988 19857 12990 19859 nw
tri 13016 19857 13018 19859 se
rect 13018 19857 13137 19859
tri 2025 19831 2051 19857 ne
rect 2051 19831 12962 19857
tri 12962 19831 12988 19857 nw
tri 12990 19831 13016 19857 se
rect 13016 19831 13137 19857
rect 1809 19803 2023 19831
tri 2023 19803 2051 19831 sw
tri 2051 19829 2053 19831 ne
rect 2053 19829 12960 19831
tri 12960 19829 12962 19831 nw
tri 12988 19829 12990 19831 se
rect 12990 19829 13137 19831
tri 2053 19803 2079 19829 ne
rect 2079 19803 12934 19829
tri 12934 19803 12960 19829 nw
tri 12962 19803 12988 19829 se
rect 12988 19803 13137 19829
rect 1809 19775 2051 19803
tri 2051 19775 2079 19803 sw
tri 2079 19801 2081 19803 ne
rect 2081 19801 12932 19803
tri 12932 19801 12934 19803 nw
tri 12960 19801 12962 19803 se
rect 12962 19801 13137 19803
tri 2081 19775 2107 19801 ne
rect 2107 19775 12906 19801
tri 12906 19775 12932 19801 nw
tri 12934 19775 12960 19801 se
rect 12960 19775 13137 19801
rect 1809 19747 2079 19775
tri 2079 19747 2107 19775 sw
tri 2107 19773 2109 19775 ne
rect 2109 19773 12904 19775
tri 12904 19773 12906 19775 nw
tri 12932 19773 12934 19775 se
rect 12934 19773 13137 19775
tri 2109 19747 2135 19773 ne
rect 2135 19747 12878 19773
tri 12878 19747 12904 19773 nw
tri 12906 19747 12932 19773 se
rect 12932 19747 13137 19773
rect 1809 19719 2107 19747
tri 2107 19719 2135 19747 sw
tri 2135 19745 2137 19747 ne
rect 2137 19745 12876 19747
tri 12876 19745 12878 19747 nw
tri 12904 19745 12906 19747 se
rect 12906 19745 13137 19747
tri 2137 19719 2163 19745 ne
rect 2163 19719 12850 19745
tri 12850 19719 12876 19745 nw
tri 12878 19719 12904 19745 se
rect 12904 19719 13137 19745
rect 1809 19697 2135 19719
rect 1566 19691 2135 19697
tri 2135 19691 2163 19719 sw
tri 2163 19717 2165 19719 ne
rect 2165 19717 12848 19719
tri 12848 19717 12850 19719 nw
tri 12876 19717 12878 19719 se
rect 12878 19717 13137 19719
tri 2165 19691 2191 19717 ne
rect 2191 19691 12822 19717
tri 12822 19691 12848 19717 nw
tri 12850 19691 12876 19717 se
rect 12876 19691 13137 19717
tri 1566 19663 1594 19691 ne
rect 1594 19663 2163 19691
tri 2163 19663 2191 19691 sw
tri 2191 19689 2193 19691 ne
rect 2193 19689 12820 19691
tri 12820 19689 12822 19691 nw
tri 12848 19689 12850 19691 se
rect 12850 19689 13137 19691
tri 2193 19663 2219 19689 ne
rect 2219 19663 12794 19689
tri 12794 19663 12820 19689 nw
tri 12822 19663 12848 19689 se
rect 12848 19663 13137 19689
tri 1594 19635 1622 19663 ne
rect 1622 19635 2191 19663
tri 2191 19635 2219 19663 sw
tri 2219 19661 2221 19663 ne
rect 2221 19661 12792 19663
tri 12792 19661 12794 19663 nw
tri 12820 19661 12822 19663 se
rect 12822 19661 13137 19663
tri 2221 19635 2247 19661 ne
rect 2247 19635 12766 19661
tri 12766 19635 12792 19661 nw
tri 12794 19635 12820 19661 se
rect 12820 19643 13137 19661
rect 13373 19857 13600 19879
tri 13600 19857 13628 19885 nw
rect 13373 19829 13572 19857
tri 13572 19829 13600 19857 nw
rect 13373 19801 13544 19829
tri 13544 19801 13572 19829 nw
rect 13373 19773 13516 19801
tri 13516 19773 13544 19801 nw
rect 13373 19745 13488 19773
tri 13488 19745 13516 19773 nw
rect 13373 19717 13460 19745
tri 13460 19717 13488 19745 nw
rect 13373 19689 13432 19717
tri 13432 19689 13460 19717 nw
rect 13373 19661 13404 19689
tri 13404 19661 13432 19689 nw
rect 13373 19643 13376 19661
rect 12820 19635 13376 19643
tri 1622 19607 1650 19635 ne
rect 1650 19613 2219 19635
rect 1650 19607 1893 19613
tri 1650 19579 1678 19607 ne
rect 1678 19579 1893 19607
tri 1678 19377 1880 19579 ne
rect 1880 19377 1893 19579
rect 2129 19607 2219 19613
tri 2219 19607 2247 19635 sw
tri 2247 19633 2249 19635 ne
rect 2249 19633 12764 19635
tri 12764 19633 12766 19635 nw
tri 12792 19633 12794 19635 se
rect 12794 19633 13376 19635
tri 13376 19633 13404 19661 nw
tri 2249 19607 2275 19633 ne
rect 2275 19607 12738 19633
tri 12738 19607 12764 19633 nw
tri 12766 19607 12792 19633 se
rect 12792 19607 13348 19633
rect 2129 19579 2247 19607
tri 2247 19579 2275 19607 sw
tri 2275 19605 2277 19607 ne
rect 2277 19605 12736 19607
tri 12736 19605 12738 19607 nw
tri 12764 19605 12766 19607 se
rect 12766 19605 13348 19607
tri 13348 19605 13376 19633 nw
tri 2277 19579 2303 19605 ne
rect 2303 19579 12710 19605
tri 12710 19579 12736 19605 nw
tri 12738 19579 12764 19605 se
rect 12764 19579 13320 19605
rect 2129 19551 2275 19579
tri 2275 19551 2303 19579 sw
tri 2303 19577 2305 19579 ne
rect 2305 19577 12708 19579
tri 12708 19577 12710 19579 nw
tri 12736 19577 12738 19579 se
rect 12738 19577 13320 19579
tri 13320 19577 13348 19605 nw
tri 2305 19551 2331 19577 ne
rect 2331 19551 12682 19577
tri 12682 19551 12708 19577 nw
tri 12710 19551 12736 19577 se
rect 12736 19559 13292 19577
rect 12736 19551 12817 19559
rect 2129 19523 2303 19551
tri 2303 19523 2331 19551 sw
tri 2331 19549 2333 19551 ne
rect 2333 19549 12680 19551
tri 12680 19549 12682 19551 nw
tri 12708 19549 12710 19551 se
rect 12710 19549 12817 19551
tri 2333 19523 2359 19549 ne
rect 2359 19523 12654 19549
tri 12654 19523 12680 19549 nw
tri 12682 19523 12708 19549 se
rect 12708 19523 12817 19549
rect 2129 19495 2331 19523
tri 2331 19495 2359 19523 sw
tri 2359 19521 2361 19523 ne
rect 2361 19521 12652 19523
tri 12652 19521 12654 19523 nw
tri 12680 19521 12682 19523 se
rect 12682 19521 12817 19523
tri 2361 19495 2387 19521 ne
rect 2387 19495 12626 19521
tri 12626 19495 12652 19521 nw
tri 12654 19495 12680 19521 se
rect 12680 19495 12817 19521
rect 2129 19467 2359 19495
tri 2359 19467 2387 19495 sw
tri 2387 19493 2389 19495 ne
rect 2389 19493 12624 19495
tri 12624 19493 12626 19495 nw
tri 12652 19493 12654 19495 se
rect 12654 19493 12817 19495
tri 2389 19467 2415 19493 ne
rect 2415 19467 12598 19493
tri 12598 19467 12624 19493 nw
tri 12626 19467 12652 19493 se
rect 12652 19467 12817 19493
rect 2129 19439 2387 19467
tri 2387 19439 2415 19467 sw
tri 2415 19465 2417 19467 ne
rect 2417 19465 12596 19467
tri 12596 19465 12598 19467 nw
tri 12624 19465 12626 19467 se
rect 12626 19465 12817 19467
tri 2417 19439 2443 19465 ne
rect 2443 19439 12570 19465
tri 12570 19439 12596 19465 nw
tri 12598 19439 12624 19465 se
rect 12624 19439 12817 19465
rect 2129 19411 2415 19439
tri 2415 19411 2443 19439 sw
tri 2443 19437 2445 19439 ne
rect 2445 19437 12568 19439
tri 12568 19437 12570 19439 nw
tri 12596 19437 12598 19439 se
rect 12598 19437 12817 19439
tri 2445 19411 2471 19437 ne
rect 2471 19411 12542 19437
tri 12542 19411 12568 19437 nw
tri 12570 19411 12596 19437 se
rect 12596 19411 12817 19437
rect 2129 19383 2443 19411
tri 2443 19383 2471 19411 sw
tri 2471 19409 2473 19411 ne
rect 2473 19409 12540 19411
tri 12540 19409 12542 19411 nw
tri 12568 19409 12570 19411 se
rect 12570 19409 12817 19411
tri 2473 19383 2499 19409 ne
rect 2499 19383 12514 19409
tri 12514 19383 12540 19409 nw
tri 12542 19383 12568 19409 se
rect 12568 19383 12817 19409
rect 2129 19377 2471 19383
tri 1880 19251 2006 19377 ne
rect 2006 19355 2471 19377
tri 2471 19355 2499 19383 sw
tri 2499 19381 2501 19383 ne
rect 2501 19381 12512 19383
tri 12512 19381 12514 19383 nw
tri 12540 19381 12542 19383 se
rect 12542 19381 12817 19383
tri 2501 19355 2527 19381 ne
rect 2527 19355 12486 19381
tri 12486 19355 12512 19381 nw
tri 12514 19355 12540 19381 se
rect 12540 19355 12817 19381
rect 2006 19335 2499 19355
tri 2499 19335 2519 19355 sw
tri 12494 19335 12514 19355 se
rect 12514 19335 12817 19355
rect 2006 19323 12817 19335
rect 13053 19549 13292 19559
tri 13292 19549 13320 19577 nw
rect 13053 19323 13066 19549
tri 13066 19323 13292 19549 nw
rect 2006 19251 12734 19323
tri 2006 19015 2242 19251 ne
rect 2242 19015 2255 19251
rect 2491 19015 2575 19251
rect 2811 19015 2895 19251
rect 3131 19015 3215 19251
rect 3451 19015 3535 19251
rect 3771 19015 3855 19251
rect 4091 19015 4175 19251
rect 4411 19015 4495 19251
rect 4731 19015 4815 19251
rect 5051 19015 5135 19251
rect 5371 19015 5455 19251
rect 5691 19015 5775 19251
rect 6011 19015 6095 19251
rect 6331 19015 6415 19251
rect 6651 19015 6735 19251
rect 6971 19015 7055 19251
rect 7291 19015 7375 19251
rect 7611 19015 7695 19251
rect 7931 19015 8015 19251
rect 8251 19015 8335 19251
rect 8571 19015 8655 19251
rect 8891 19015 8975 19251
rect 9211 19015 9295 19251
rect 9531 19015 9615 19251
rect 9851 19015 9935 19251
rect 10171 19015 10255 19251
rect 10491 19015 10575 19251
rect 10811 19015 10895 19251
rect 11131 19015 11215 19251
rect 11451 19015 11535 19251
rect 11771 19015 11855 19251
rect 12091 19015 12175 19251
rect 12411 19015 12495 19251
rect 12731 19015 12734 19251
tri 2242 18991 2266 19015 ne
rect 2266 18991 12734 19015
tri 12734 18991 13066 19323 nw
<< rm5 >>
tri 2405 33663 2425 33683 se
rect 2425 33663 12578 33683
tri 12578 33663 12598 33683 sw
tri 2390 33648 2405 33663 se
rect 2405 33648 2418 33663
tri 2418 33648 2433 33663 nw
tri 12570 33648 12585 33663 ne
rect 12585 33648 12598 33663
tri 12598 33648 12613 33663 sw
tri 2362 33620 2390 33648 se
rect 2390 33635 2405 33648
tri 2405 33635 2418 33648 nw
tri 12585 33635 12598 33648 ne
rect 12598 33635 12613 33648
tri 12613 33635 12626 33648 sw
tri 2390 33620 2405 33635 nw
tri 12598 33620 12613 33635 ne
rect 12613 33620 12626 33635
tri 12626 33620 12641 33635 sw
tri 2334 33592 2362 33620 se
rect 2362 33607 2377 33620
tri 2377 33607 2390 33620 nw
tri 12613 33607 12626 33620 ne
rect 12626 33607 12641 33620
tri 12641 33607 12654 33620 sw
tri 2362 33592 2377 33607 nw
tri 12626 33592 12641 33607 ne
rect 12641 33592 12654 33607
tri 12654 33592 12669 33607 sw
tri 2306 33564 2334 33592 se
rect 2334 33579 2349 33592
tri 2349 33579 2362 33592 nw
tri 12641 33579 12654 33592 ne
rect 12654 33579 12669 33592
tri 12669 33579 12682 33592 sw
tri 2334 33564 2349 33579 nw
tri 12654 33564 12669 33579 ne
rect 12669 33564 12682 33579
tri 12682 33564 12697 33579 sw
tri 2278 33536 2306 33564 se
rect 2306 33551 2321 33564
tri 2321 33551 2334 33564 nw
tri 12669 33551 12682 33564 ne
rect 12682 33551 12697 33564
tri 12697 33551 12710 33564 sw
tri 2306 33536 2321 33551 nw
tri 12682 33536 12697 33551 ne
rect 12697 33536 12710 33551
tri 12710 33536 12725 33551 sw
tri 2250 33508 2278 33536 se
rect 2278 33523 2293 33536
tri 2293 33523 2306 33536 nw
tri 12697 33523 12710 33536 ne
rect 12710 33523 12725 33536
tri 12725 33523 12738 33536 sw
tri 2278 33508 2293 33523 nw
tri 12710 33508 12725 33523 ne
rect 12725 33508 12738 33523
tri 12738 33508 12753 33523 sw
tri 2222 33480 2250 33508 se
rect 2250 33495 2265 33508
tri 2265 33495 2278 33508 nw
tri 12725 33495 12738 33508 ne
rect 12738 33495 12753 33508
tri 12753 33495 12766 33508 sw
tri 2250 33480 2265 33495 nw
tri 12738 33480 12753 33495 ne
rect 12753 33480 12766 33495
tri 12766 33480 12781 33495 sw
tri 2194 33452 2222 33480 se
rect 2222 33467 2237 33480
tri 2237 33467 2250 33480 nw
tri 12753 33467 12766 33480 ne
rect 12766 33467 12781 33480
tri 12781 33467 12794 33480 sw
tri 2222 33452 2237 33467 nw
tri 12766 33452 12781 33467 ne
rect 12781 33452 12794 33467
tri 12794 33452 12809 33467 sw
tri 2166 33424 2194 33452 se
rect 2194 33439 2209 33452
tri 2209 33439 2222 33452 nw
tri 12781 33439 12794 33452 ne
rect 12794 33439 12809 33452
tri 12809 33439 12822 33452 sw
tri 2194 33424 2209 33439 nw
tri 12794 33424 12809 33439 ne
rect 12809 33424 12822 33439
tri 12822 33424 12837 33439 sw
tri 2138 33396 2166 33424 se
rect 2166 33411 2181 33424
tri 2181 33411 2194 33424 nw
tri 12809 33411 12822 33424 ne
rect 12822 33411 12837 33424
tri 12837 33411 12850 33424 sw
tri 2166 33396 2181 33411 nw
tri 12822 33396 12837 33411 ne
rect 12837 33396 12850 33411
tri 12850 33396 12865 33411 sw
tri 2110 33368 2138 33396 se
rect 2138 33383 2153 33396
tri 2153 33383 2166 33396 nw
tri 12837 33383 12850 33396 ne
rect 12850 33383 12865 33396
tri 12865 33383 12878 33396 sw
tri 2138 33368 2153 33383 nw
tri 12850 33368 12865 33383 ne
rect 12865 33368 12878 33383
tri 12878 33368 12893 33383 sw
tri 2082 33340 2110 33368 se
rect 2110 33355 2125 33368
tri 2125 33355 2138 33368 nw
tri 12865 33355 12878 33368 ne
rect 12878 33355 12893 33368
tri 12893 33355 12906 33368 sw
tri 2110 33340 2125 33355 nw
tri 12878 33340 12893 33355 ne
rect 12893 33340 12906 33355
tri 12906 33340 12921 33355 sw
tri 2054 33312 2082 33340 se
rect 2082 33327 2097 33340
tri 2097 33327 2110 33340 nw
tri 12893 33327 12906 33340 ne
rect 12906 33327 12921 33340
tri 12921 33327 12934 33340 sw
tri 2082 33312 2097 33327 nw
tri 12906 33312 12921 33327 ne
rect 12921 33312 12934 33327
tri 12934 33312 12949 33327 sw
tri 2026 33284 2054 33312 se
rect 2054 33299 2069 33312
tri 2069 33299 2082 33312 nw
tri 12921 33299 12934 33312 ne
rect 12934 33299 12949 33312
tri 12949 33299 12962 33312 sw
tri 2054 33284 2069 33299 nw
tri 12934 33284 12949 33299 ne
rect 12949 33284 12962 33299
tri 12962 33284 12977 33299 sw
tri 1998 33256 2026 33284 se
rect 2026 33271 2041 33284
tri 2041 33271 2054 33284 nw
tri 12949 33271 12962 33284 ne
rect 12962 33271 12977 33284
tri 12977 33271 12990 33284 sw
tri 2026 33256 2041 33271 nw
tri 12962 33256 12977 33271 ne
rect 12977 33256 12990 33271
tri 12990 33256 13005 33271 sw
tri 1970 33228 1998 33256 se
rect 1998 33243 2013 33256
tri 2013 33243 2026 33256 nw
tri 12977 33243 12990 33256 ne
rect 12990 33243 13005 33256
tri 13005 33243 13018 33256 sw
tri 1998 33228 2013 33243 nw
tri 12990 33228 13005 33243 ne
rect 13005 33228 13018 33243
tri 13018 33228 13033 33243 sw
tri 1942 33200 1970 33228 se
rect 1970 33215 1985 33228
tri 1985 33215 1998 33228 nw
tri 13005 33215 13018 33228 ne
rect 13018 33215 13033 33228
tri 13033 33215 13046 33228 sw
tri 1970 33200 1985 33215 nw
tri 13018 33200 13033 33215 ne
rect 13033 33200 13046 33215
tri 13046 33200 13061 33215 sw
tri 1914 33172 1942 33200 se
rect 1942 33187 1957 33200
tri 1957 33187 1970 33200 nw
tri 13033 33187 13046 33200 ne
rect 13046 33187 13061 33200
tri 13061 33187 13074 33200 sw
tri 1942 33172 1957 33187 nw
tri 13046 33172 13061 33187 ne
rect 13061 33172 13074 33187
tri 13074 33172 13089 33187 sw
tri 1886 33144 1914 33172 se
rect 1914 33159 1929 33172
tri 1929 33159 1942 33172 nw
tri 13061 33159 13074 33172 ne
rect 13074 33159 13089 33172
tri 13089 33159 13102 33172 sw
tri 1914 33144 1929 33159 nw
tri 13074 33144 13089 33159 ne
rect 13089 33144 13102 33159
tri 13102 33144 13117 33159 sw
tri 1858 33116 1886 33144 se
rect 1886 33131 1901 33144
tri 1901 33131 1914 33144 nw
tri 13089 33131 13102 33144 ne
rect 13102 33131 13117 33144
tri 13117 33131 13130 33144 sw
tri 1886 33116 1901 33131 nw
tri 13102 33116 13117 33131 ne
rect 13117 33116 13130 33131
tri 13130 33116 13145 33131 sw
tri 1830 33088 1858 33116 se
rect 1858 33103 1873 33116
tri 1873 33103 1886 33116 nw
tri 13117 33103 13130 33116 ne
rect 13130 33103 13145 33116
tri 13145 33103 13158 33116 sw
tri 1858 33088 1873 33103 nw
tri 13130 33088 13145 33103 ne
rect 13145 33088 13158 33103
tri 13158 33088 13173 33103 sw
tri 1802 33060 1830 33088 se
rect 1830 33075 1845 33088
tri 1845 33075 1858 33088 nw
tri 13145 33075 13158 33088 ne
rect 13158 33075 13173 33088
tri 13173 33075 13186 33088 sw
tri 1830 33060 1845 33075 nw
tri 13158 33060 13173 33075 ne
rect 13173 33060 13186 33075
tri 13186 33060 13201 33075 sw
tri 1774 33032 1802 33060 se
rect 1802 33047 1817 33060
tri 1817 33047 1830 33060 nw
tri 13173 33047 13186 33060 ne
rect 13186 33047 13201 33060
tri 13201 33047 13214 33060 sw
tri 1802 33032 1817 33047 nw
tri 13186 33032 13201 33047 ne
rect 13201 33032 13214 33047
tri 13214 33032 13229 33047 sw
tri 1746 33004 1774 33032 se
rect 1774 33019 1789 33032
tri 1789 33019 1802 33032 nw
tri 13201 33019 13214 33032 ne
rect 13214 33019 13229 33032
tri 13229 33019 13242 33032 sw
tri 1774 33004 1789 33019 nw
tri 13214 33004 13229 33019 ne
rect 13229 33004 13242 33019
tri 13242 33004 13257 33019 sw
tri 1718 32976 1746 33004 se
rect 1746 32991 1761 33004
tri 1761 32991 1774 33004 nw
tri 13229 32991 13242 33004 ne
rect 13242 32991 13257 33004
tri 13257 32991 13270 33004 sw
tri 1746 32976 1761 32991 nw
tri 13242 32976 13257 32991 ne
rect 13257 32976 13270 32991
tri 13270 32976 13285 32991 sw
tri 1690 32948 1718 32976 se
rect 1718 32963 1733 32976
tri 1733 32963 1746 32976 nw
tri 13257 32963 13270 32976 ne
rect 13270 32963 13285 32976
tri 13285 32963 13298 32976 sw
tri 1718 32948 1733 32963 nw
tri 13270 32948 13285 32963 ne
rect 13285 32948 13298 32963
tri 13298 32948 13313 32963 sw
tri 1662 32920 1690 32948 se
rect 1690 32935 1705 32948
tri 1705 32935 1718 32948 nw
tri 13285 32935 13298 32948 ne
rect 13298 32935 13313 32948
tri 13313 32935 13326 32948 sw
tri 1690 32920 1705 32935 nw
tri 13298 32920 13313 32935 ne
rect 13313 32920 13326 32935
tri 13326 32920 13341 32935 sw
tri 1634 32892 1662 32920 se
rect 1662 32907 1677 32920
tri 1677 32907 1690 32920 nw
tri 13313 32907 13326 32920 ne
rect 13326 32907 13341 32920
tri 13341 32907 13354 32920 sw
tri 1662 32892 1677 32907 nw
tri 13326 32892 13341 32907 ne
rect 13341 32892 13354 32907
tri 13354 32892 13369 32907 sw
tri 1606 32864 1634 32892 se
rect 1634 32879 1649 32892
tri 1649 32879 1662 32892 nw
tri 13341 32879 13354 32892 ne
rect 13354 32879 13369 32892
tri 13369 32879 13382 32892 sw
tri 1634 32864 1649 32879 nw
tri 13354 32864 13369 32879 ne
rect 13369 32864 13382 32879
tri 13382 32864 13397 32879 sw
tri 1578 32836 1606 32864 se
rect 1606 32851 1621 32864
tri 1621 32851 1634 32864 nw
tri 13369 32851 13382 32864 ne
rect 13382 32851 13397 32864
tri 13397 32851 13410 32864 sw
tri 1606 32836 1621 32851 nw
tri 13382 32836 13397 32851 ne
rect 13397 32836 13410 32851
tri 13410 32836 13425 32851 sw
tri 1550 32808 1578 32836 se
rect 1578 32823 1593 32836
tri 1593 32823 1606 32836 nw
tri 13397 32823 13410 32836 ne
rect 13410 32823 13425 32836
tri 13425 32823 13438 32836 sw
tri 1578 32808 1593 32823 nw
tri 13410 32808 13425 32823 ne
rect 13425 32808 13438 32823
tri 13438 32808 13453 32823 sw
tri 1522 32780 1550 32808 se
rect 1550 32795 1565 32808
tri 1565 32795 1578 32808 nw
tri 13425 32795 13438 32808 ne
rect 13438 32795 13453 32808
tri 13453 32795 13466 32808 sw
tri 1550 32780 1565 32795 nw
tri 13438 32780 13453 32795 ne
rect 13453 32780 13466 32795
tri 13466 32780 13481 32795 sw
tri 1507 32765 1522 32780 se
rect 1522 32767 1537 32780
tri 1537 32767 1550 32780 nw
tri 13453 32767 13466 32780 ne
rect 13466 32767 13481 32780
tri 13481 32767 13494 32780 sw
rect 1522 32765 1535 32767
tri 1535 32765 1537 32767 nw
tri 13466 32765 13468 32767 ne
rect 13468 32765 13494 32767
tri 13494 32765 13496 32767 sw
tri 1494 32752 1507 32765 se
rect 1507 32752 1522 32765
tri 1522 32752 1535 32765 nw
tri 13468 32752 13481 32765 ne
rect 13481 32752 13496 32765
tri 13496 32752 13509 32765 sw
tri 1466 32724 1494 32752 se
rect 1494 32739 1509 32752
tri 1509 32739 1522 32752 nw
tri 13481 32739 13494 32752 ne
rect 13494 32739 13509 32752
tri 13509 32739 13522 32752 sw
tri 1494 32724 1509 32739 nw
tri 13494 32724 13509 32739 ne
rect 13509 32724 13522 32739
tri 13522 32724 13537 32739 sw
tri 1438 32696 1466 32724 se
rect 1466 32711 1481 32724
tri 1481 32711 1494 32724 nw
tri 13509 32711 13522 32724 ne
rect 13522 32711 13537 32724
tri 13537 32711 13550 32724 sw
tri 1466 32696 1481 32711 nw
tri 13522 32696 13537 32711 ne
rect 13537 32696 13550 32711
tri 13550 32696 13565 32711 sw
tri 1410 32668 1438 32696 se
rect 1438 32683 1453 32696
tri 1453 32683 1466 32696 nw
tri 13537 32683 13550 32696 ne
rect 13550 32683 13565 32696
tri 13565 32683 13578 32696 sw
tri 1438 32668 1453 32683 nw
tri 13550 32668 13565 32683 ne
rect 13565 32668 13578 32683
tri 13578 32668 13593 32683 sw
tri 1382 32640 1410 32668 se
rect 1410 32655 1425 32668
tri 1425 32655 1438 32668 nw
tri 13565 32655 13578 32668 ne
rect 13578 32657 13593 32668
tri 13593 32657 13604 32668 sw
rect 13578 32655 13604 32657
tri 13604 32655 13606 32657 sw
tri 1410 32640 1425 32655 nw
tri 13578 32640 13593 32655 ne
rect 13593 32640 13606 32655
tri 13606 32640 13621 32655 sw
tri 1354 32612 1382 32640 se
rect 1382 32629 1399 32640
tri 1399 32629 1410 32640 nw
tri 13593 32629 13604 32640 ne
rect 13604 32637 13621 32640
tri 13621 32637 13624 32640 sw
tri 1382 32612 1399 32629 nw
tri 1334 32592 1354 32612 se
rect 1354 32592 1362 32612
tri 1362 32592 1382 32612 nw
rect 1334 20520 1354 32592
tri 1354 32584 1362 32592 nw
tri 1354 20520 1362 20528 sw
tri 1334 20503 1351 20520 ne
rect 1351 20503 1362 20520
tri 1362 20503 1379 20520 sw
tri 1351 20500 1354 20503 ne
rect 1354 20500 1379 20503
tri 1379 20500 1382 20503 sw
tri 1354 20475 1379 20500 ne
rect 1379 20475 1382 20500
tri 1382 20475 1407 20500 sw
tri 1379 20447 1407 20475 ne
tri 1407 20473 1409 20475 sw
rect 1407 20447 1409 20473
tri 1409 20447 1435 20473 sw
tri 13578 20447 13604 20473 se
rect 13604 20465 13624 32637
rect 13604 20447 13606 20465
tri 13606 20447 13624 20465 nw
tri 1407 20419 1435 20447 ne
tri 1435 20445 1437 20447 sw
tri 13576 20445 13578 20447 se
rect 13578 20445 13604 20447
tri 13604 20445 13606 20447 nw
rect 1435 20419 1437 20445
tri 1437 20419 1463 20445 sw
tri 13550 20419 13576 20445 se
rect 13576 20419 13578 20445
tri 13578 20419 13604 20445 nw
tri 1435 20391 1463 20419 ne
tri 1463 20417 1465 20419 sw
tri 13548 20417 13550 20419 se
rect 13550 20417 13576 20419
tri 13576 20417 13578 20419 nw
rect 1463 20391 1465 20417
tri 1465 20391 1491 20417 sw
tri 13522 20391 13548 20417 se
rect 13548 20391 13550 20417
tri 13550 20391 13576 20417 nw
tri 1463 20363 1491 20391 ne
tri 1491 20389 1493 20391 sw
tri 13520 20389 13522 20391 se
rect 13522 20389 13548 20391
tri 13548 20389 13550 20391 nw
rect 1491 20363 1493 20389
tri 1493 20363 1519 20389 sw
tri 13494 20363 13520 20389 se
rect 13520 20363 13522 20389
tri 13522 20363 13548 20389 nw
tri 1491 20335 1519 20363 ne
tri 1519 20361 1521 20363 sw
tri 13492 20361 13494 20363 se
rect 13494 20361 13520 20363
tri 13520 20361 13522 20363 nw
rect 1519 20335 1521 20361
tri 1521 20335 1547 20361 sw
tri 13466 20335 13492 20361 se
rect 13492 20335 13494 20361
tri 13494 20335 13520 20361 nw
tri 1519 20307 1547 20335 ne
tri 1547 20333 1549 20335 sw
tri 13464 20333 13466 20335 se
rect 13466 20333 13492 20335
tri 13492 20333 13494 20335 nw
rect 1547 20307 1549 20333
tri 1549 20307 1575 20333 sw
tri 13438 20307 13464 20333 se
rect 13464 20307 13466 20333
tri 13466 20307 13492 20333 nw
tri 1547 20297 1557 20307 ne
rect 1557 20305 1575 20307
tri 1575 20305 1577 20307 sw
tri 13436 20305 13438 20307 se
rect 13438 20305 13464 20307
tri 13464 20305 13466 20307 nw
rect 1557 20297 1577 20305
tri 1577 20297 1585 20305 sw
tri 13428 20297 13436 20305 se
rect 13436 20297 13456 20305
tri 13456 20297 13464 20305 nw
tri 1557 20279 1575 20297 ne
rect 1575 20279 1585 20297
tri 1585 20279 1603 20297 sw
tri 13410 20279 13428 20297 se
rect 13428 20279 13438 20297
tri 13438 20279 13456 20297 nw
tri 1575 20251 1603 20279 ne
tri 1603 20277 1605 20279 sw
tri 13408 20277 13410 20279 se
rect 13410 20277 13436 20279
tri 13436 20277 13438 20279 nw
rect 1603 20251 1605 20277
tri 1605 20251 1631 20277 sw
tri 13382 20251 13408 20277 se
rect 13408 20251 13410 20277
tri 13410 20251 13436 20277 nw
tri 1603 20223 1631 20251 ne
tri 1631 20249 1633 20251 sw
tri 13380 20249 13382 20251 se
rect 13382 20249 13408 20251
tri 13408 20249 13410 20251 nw
rect 1631 20223 1633 20249
tri 1633 20223 1659 20249 sw
tri 13354 20223 13380 20249 se
rect 13380 20223 13382 20249
tri 13382 20223 13408 20249 nw
tri 1631 20195 1659 20223 ne
tri 1659 20221 1661 20223 sw
tri 13352 20221 13354 20223 se
rect 13354 20221 13380 20223
tri 13380 20221 13382 20223 nw
rect 1659 20195 1661 20221
tri 1661 20195 1687 20221 sw
tri 13326 20195 13352 20221 se
rect 13352 20195 13354 20221
tri 13354 20195 13380 20221 nw
tri 1659 20167 1687 20195 ne
tri 1687 20193 1689 20195 sw
tri 13324 20193 13326 20195 se
rect 13326 20193 13352 20195
tri 13352 20193 13354 20195 nw
rect 1687 20167 1689 20193
tri 1689 20167 1715 20193 sw
tri 13298 20167 13324 20193 se
rect 13324 20167 13326 20193
tri 13326 20167 13352 20193 nw
tri 1687 20139 1715 20167 ne
tri 1715 20165 1717 20167 sw
tri 13296 20165 13298 20167 se
rect 13298 20165 13324 20167
tri 13324 20165 13326 20167 nw
rect 1715 20139 1717 20165
tri 1717 20139 1743 20165 sw
tri 13270 20139 13296 20165 se
rect 13296 20139 13298 20165
tri 13298 20139 13324 20165 nw
tri 1715 20111 1743 20139 ne
tri 1743 20137 1745 20139 sw
tri 13268 20137 13270 20139 se
rect 13270 20137 13296 20139
tri 13296 20137 13298 20139 nw
rect 1743 20111 1745 20137
tri 1745 20111 1771 20137 sw
tri 13242 20111 13268 20137 se
rect 13268 20111 13270 20137
tri 13270 20111 13296 20137 nw
tri 1743 20083 1771 20111 ne
tri 1771 20109 1773 20111 sw
tri 13240 20109 13242 20111 se
rect 13242 20109 13268 20111
tri 13268 20109 13270 20111 nw
rect 1771 20083 1773 20109
tri 1773 20083 1799 20109 sw
tri 13214 20083 13240 20109 se
rect 13240 20083 13242 20109
tri 13242 20083 13268 20109 nw
tri 1771 20055 1799 20083 ne
tri 1799 20081 1801 20083 sw
tri 13212 20081 13214 20083 se
rect 13214 20081 13240 20083
tri 13240 20081 13242 20083 nw
rect 1799 20055 1801 20081
tri 1801 20055 1827 20081 sw
tri 13186 20055 13212 20081 se
rect 13212 20055 13214 20081
tri 13214 20055 13240 20081 nw
tri 1799 20027 1827 20055 ne
tri 1827 20053 1829 20055 sw
tri 13184 20053 13186 20055 se
rect 13186 20053 13212 20055
tri 13212 20053 13214 20055 nw
rect 1827 20027 1829 20053
tri 1829 20027 1855 20053 sw
tri 13158 20027 13184 20053 se
rect 13184 20027 13186 20053
tri 13186 20027 13212 20053 nw
tri 1827 19999 1855 20027 ne
tri 1855 20025 1857 20027 sw
tri 13156 20025 13158 20027 se
rect 13158 20025 13184 20027
tri 13184 20025 13186 20027 nw
rect 1855 19999 1857 20025
tri 1857 19999 1883 20025 sw
tri 13130 19999 13156 20025 se
rect 13156 19999 13158 20025
tri 13158 19999 13184 20025 nw
tri 1855 19971 1883 19999 ne
tri 1883 19997 1885 19999 sw
tri 13128 19997 13130 19999 se
rect 13130 19997 13156 19999
tri 13156 19997 13158 19999 nw
rect 1883 19971 1885 19997
tri 1885 19971 1911 19997 sw
tri 13102 19971 13128 19997 se
rect 13128 19971 13130 19997
tri 13130 19971 13156 19997 nw
tri 1883 19943 1911 19971 ne
tri 1911 19969 1913 19971 sw
tri 13100 19969 13102 19971 se
rect 13102 19969 13128 19971
tri 13128 19969 13130 19971 nw
rect 1911 19943 1913 19969
tri 1913 19943 1939 19969 sw
tri 13074 19943 13100 19969 se
rect 13100 19943 13102 19969
tri 13102 19943 13128 19969 nw
tri 1911 19915 1939 19943 ne
tri 1939 19941 1941 19943 sw
tri 13072 19941 13074 19943 se
rect 13074 19941 13100 19943
tri 13100 19941 13102 19943 nw
rect 1939 19915 1941 19941
tri 1941 19915 1967 19941 sw
tri 13046 19915 13072 19941 se
rect 13072 19915 13074 19941
tri 13074 19915 13100 19941 nw
tri 1939 19887 1967 19915 ne
tri 1967 19913 1969 19915 sw
tri 13044 19913 13046 19915 se
rect 13046 19913 13072 19915
tri 13072 19913 13074 19915 nw
rect 1967 19887 1969 19913
tri 1969 19887 1995 19913 sw
tri 13018 19887 13044 19913 se
rect 13044 19887 13046 19913
tri 13046 19887 13072 19913 nw
tri 1967 19859 1995 19887 ne
tri 1995 19885 1997 19887 sw
tri 13016 19885 13018 19887 se
rect 13018 19885 13044 19887
tri 13044 19885 13046 19887 nw
rect 1995 19859 1997 19885
tri 1997 19859 2023 19885 sw
tri 12990 19859 13016 19885 se
rect 13016 19859 13018 19885
tri 13018 19859 13044 19885 nw
tri 1995 19831 2023 19859 ne
tri 2023 19857 2025 19859 sw
tri 12988 19857 12990 19859 se
rect 12990 19857 13016 19859
tri 13016 19857 13018 19859 nw
rect 2023 19831 2025 19857
tri 2025 19831 2051 19857 sw
tri 12962 19831 12988 19857 se
rect 12988 19831 12990 19857
tri 12990 19831 13016 19857 nw
tri 2023 19803 2051 19831 ne
tri 2051 19829 2053 19831 sw
tri 12960 19829 12962 19831 se
rect 12962 19829 12988 19831
tri 12988 19829 12990 19831 nw
rect 2051 19803 2053 19829
tri 2053 19803 2079 19829 sw
tri 12934 19803 12960 19829 se
rect 12960 19803 12962 19829
tri 12962 19803 12988 19829 nw
tri 2051 19775 2079 19803 ne
tri 2079 19801 2081 19803 sw
tri 12932 19801 12934 19803 se
rect 12934 19801 12960 19803
tri 12960 19801 12962 19803 nw
rect 2079 19775 2081 19801
tri 2081 19775 2107 19801 sw
tri 12906 19775 12932 19801 se
rect 12932 19775 12934 19801
tri 12934 19775 12960 19801 nw
tri 2079 19747 2107 19775 ne
tri 2107 19773 2109 19775 sw
tri 12904 19773 12906 19775 se
rect 12906 19773 12932 19775
tri 12932 19773 12934 19775 nw
rect 2107 19747 2109 19773
tri 2109 19747 2135 19773 sw
tri 12878 19747 12904 19773 se
rect 12904 19747 12906 19773
tri 12906 19747 12932 19773 nw
tri 2107 19719 2135 19747 ne
tri 2135 19745 2137 19747 sw
tri 12876 19745 12878 19747 se
rect 12878 19745 12904 19747
tri 12904 19745 12906 19747 nw
rect 2135 19719 2137 19745
tri 2137 19719 2163 19745 sw
tri 12850 19719 12876 19745 se
rect 12876 19719 12878 19745
tri 12878 19719 12904 19745 nw
tri 2135 19691 2163 19719 ne
tri 2163 19717 2165 19719 sw
tri 12848 19717 12850 19719 se
rect 12850 19717 12876 19719
tri 12876 19717 12878 19719 nw
rect 2163 19691 2165 19717
tri 2165 19691 2191 19717 sw
tri 12822 19691 12848 19717 se
rect 12848 19691 12850 19717
tri 12850 19691 12876 19717 nw
tri 2163 19663 2191 19691 ne
tri 2191 19689 2193 19691 sw
tri 12820 19689 12822 19691 se
rect 12822 19689 12848 19691
tri 12848 19689 12850 19691 nw
rect 2191 19663 2193 19689
tri 2193 19663 2219 19689 sw
tri 12794 19663 12820 19689 se
rect 12820 19663 12822 19689
tri 12822 19663 12848 19689 nw
tri 2191 19635 2219 19663 ne
tri 2219 19661 2221 19663 sw
tri 12792 19661 12794 19663 se
rect 12794 19661 12820 19663
tri 12820 19661 12822 19663 nw
rect 2219 19635 2221 19661
tri 2221 19635 2247 19661 sw
tri 12766 19635 12792 19661 se
rect 12792 19635 12794 19661
tri 12794 19635 12820 19661 nw
tri 2219 19607 2247 19635 ne
tri 2247 19633 2249 19635 sw
tri 12764 19633 12766 19635 se
rect 12766 19633 12792 19635
tri 12792 19633 12794 19635 nw
rect 2247 19607 2249 19633
tri 2249 19607 2275 19633 sw
tri 12738 19607 12764 19633 se
rect 12764 19607 12766 19633
tri 12766 19607 12792 19633 nw
tri 2247 19579 2275 19607 ne
tri 2275 19605 2277 19607 sw
tri 12736 19605 12738 19607 se
rect 12738 19605 12764 19607
tri 12764 19605 12766 19607 nw
rect 2275 19579 2277 19605
tri 2277 19579 2303 19605 sw
tri 12710 19579 12736 19605 se
rect 12736 19579 12738 19605
tri 12738 19579 12764 19605 nw
tri 2275 19551 2303 19579 ne
tri 2303 19577 2305 19579 sw
tri 12708 19577 12710 19579 se
rect 12710 19577 12736 19579
tri 12736 19577 12738 19579 nw
rect 2303 19551 2305 19577
tri 2305 19551 2331 19577 sw
tri 12682 19551 12708 19577 se
rect 12708 19551 12710 19577
tri 12710 19551 12736 19577 nw
tri 2303 19523 2331 19551 ne
tri 2331 19549 2333 19551 sw
tri 12680 19549 12682 19551 se
rect 12682 19549 12708 19551
tri 12708 19549 12710 19551 nw
rect 2331 19523 2333 19549
tri 2333 19523 2359 19549 sw
tri 12654 19523 12680 19549 se
rect 12680 19523 12682 19549
tri 12682 19523 12708 19549 nw
tri 2331 19495 2359 19523 ne
tri 2359 19521 2361 19523 sw
tri 12652 19521 12654 19523 se
rect 12654 19521 12680 19523
tri 12680 19521 12682 19523 nw
rect 2359 19495 2361 19521
tri 2361 19495 2387 19521 sw
tri 12626 19495 12652 19521 se
rect 12652 19495 12654 19521
tri 12654 19495 12680 19521 nw
tri 2359 19467 2387 19495 ne
tri 2387 19493 2389 19495 sw
tri 12624 19493 12626 19495 se
rect 12626 19493 12652 19495
tri 12652 19493 12654 19495 nw
rect 2387 19467 2389 19493
tri 2389 19467 2415 19493 sw
tri 12598 19467 12624 19493 se
rect 12624 19467 12626 19493
tri 12626 19467 12652 19493 nw
tri 2387 19439 2415 19467 ne
tri 2415 19465 2417 19467 sw
tri 12596 19465 12598 19467 se
rect 12598 19465 12624 19467
tri 12624 19465 12626 19467 nw
rect 2415 19439 2417 19465
tri 2417 19439 2443 19465 sw
tri 12570 19439 12596 19465 se
rect 12596 19439 12598 19465
tri 12598 19439 12624 19465 nw
tri 2415 19411 2443 19439 ne
tri 2443 19437 2445 19439 sw
tri 12568 19437 12570 19439 se
rect 12570 19437 12596 19439
tri 12596 19437 12598 19439 nw
rect 2443 19411 2445 19437
tri 2445 19411 2471 19437 sw
tri 12542 19411 12568 19437 se
rect 12568 19411 12570 19437
tri 12570 19411 12596 19437 nw
tri 2443 19383 2471 19411 ne
tri 2471 19409 2473 19411 sw
tri 12540 19409 12542 19411 se
rect 12542 19409 12568 19411
tri 12568 19409 12570 19411 nw
rect 2471 19383 2473 19409
tri 2473 19383 2499 19409 sw
tri 12514 19383 12540 19409 se
rect 12540 19383 12542 19409
tri 12542 19383 12568 19409 nw
tri 2471 19355 2499 19383 ne
tri 2499 19381 2501 19383 sw
tri 12512 19381 12514 19383 se
rect 12514 19381 12540 19383
tri 12540 19381 12542 19383 nw
rect 2499 19355 2501 19381
tri 2501 19355 2527 19381 sw
tri 12486 19355 12512 19381 se
rect 12512 19355 12514 19381
tri 12514 19355 12540 19381 nw
tri 2499 19335 2519 19355 ne
rect 2519 19335 12494 19355
tri 12494 19335 12514 19355 nw
<< glass >>
tri 1500 32541 2490 33531 se
rect 2490 32541 12510 33531
tri 12510 32541 13500 33531 sw
rect 1500 20521 13500 32541
tri 1500 19531 2490 20521 ne
rect 2490 19531 12510 20521
tri 12510 19531 13500 20521 nw
use sky130_fd_pr__padplhp__example_559591418080  sky130_fd_pr__padplhp__example_559591418080_0
timestamp 1676037725
transform 1 0 1500 0 1 19531
box -478 -478 1 1
<< properties >>
string GDS_END 8190624
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8190360
<< end >>
